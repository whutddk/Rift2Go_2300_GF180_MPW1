magic
tech gf180mcuD
magscale 1 5
timestamp 1698895503
<< obsm1 >>
rect 672 855 286328 287265
<< metal2 >>
rect 4256 288439 4312 288839
rect 12208 288439 12264 288839
rect 20160 288439 20216 288839
rect 28112 288439 28168 288839
rect 36064 288439 36120 288839
rect 44016 288439 44072 288839
rect 51968 288439 52024 288839
rect 59920 288439 59976 288839
rect 67872 288439 67928 288839
rect 75824 288439 75880 288839
rect 83776 288439 83832 288839
rect 91728 288439 91784 288839
rect 99680 288439 99736 288839
rect 107632 288439 107688 288839
rect 115584 288439 115640 288839
rect 123536 288439 123592 288839
rect 131488 288439 131544 288839
rect 139440 288439 139496 288839
rect 147392 288439 147448 288839
rect 155344 288439 155400 288839
rect 163296 288439 163352 288839
rect 171248 288439 171304 288839
rect 179200 288439 179256 288839
rect 187152 288439 187208 288839
rect 195104 288439 195160 288839
rect 203056 288439 203112 288839
rect 211008 288439 211064 288839
rect 218960 288439 219016 288839
rect 226912 288439 226968 288839
rect 234864 288439 234920 288839
rect 242816 288439 242872 288839
rect 250768 288439 250824 288839
rect 258720 288439 258776 288839
rect 266672 288439 266728 288839
rect 274624 288439 274680 288839
rect 282576 288439 282632 288839
rect 8624 0 8680 400
rect 9520 0 9576 400
rect 10416 0 10472 400
rect 11312 0 11368 400
rect 12208 0 12264 400
rect 13104 0 13160 400
rect 14000 0 14056 400
rect 14896 0 14952 400
rect 15792 0 15848 400
rect 16688 0 16744 400
rect 17584 0 17640 400
rect 18480 0 18536 400
rect 19376 0 19432 400
rect 20272 0 20328 400
rect 21168 0 21224 400
rect 22064 0 22120 400
rect 22960 0 23016 400
rect 23856 0 23912 400
rect 24752 0 24808 400
rect 25648 0 25704 400
rect 26544 0 26600 400
rect 27440 0 27496 400
rect 28336 0 28392 400
rect 29232 0 29288 400
rect 30128 0 30184 400
rect 31024 0 31080 400
rect 31920 0 31976 400
rect 32816 0 32872 400
rect 33712 0 33768 400
rect 34608 0 34664 400
rect 35504 0 35560 400
rect 36400 0 36456 400
rect 37296 0 37352 400
rect 38192 0 38248 400
rect 39088 0 39144 400
rect 39984 0 40040 400
rect 40880 0 40936 400
rect 41776 0 41832 400
rect 42672 0 42728 400
rect 43568 0 43624 400
rect 44464 0 44520 400
rect 45360 0 45416 400
rect 46256 0 46312 400
rect 47152 0 47208 400
rect 48048 0 48104 400
rect 48944 0 49000 400
rect 49840 0 49896 400
rect 50736 0 50792 400
rect 51632 0 51688 400
rect 52528 0 52584 400
rect 53424 0 53480 400
rect 54320 0 54376 400
rect 55216 0 55272 400
rect 56112 0 56168 400
rect 57008 0 57064 400
rect 57904 0 57960 400
rect 58800 0 58856 400
rect 59696 0 59752 400
rect 60592 0 60648 400
rect 61488 0 61544 400
rect 62384 0 62440 400
rect 63280 0 63336 400
rect 64176 0 64232 400
rect 65072 0 65128 400
rect 65968 0 66024 400
rect 66864 0 66920 400
rect 67760 0 67816 400
rect 68656 0 68712 400
rect 69552 0 69608 400
rect 70448 0 70504 400
rect 71344 0 71400 400
rect 72240 0 72296 400
rect 73136 0 73192 400
rect 74032 0 74088 400
rect 74928 0 74984 400
rect 75824 0 75880 400
rect 76720 0 76776 400
rect 77616 0 77672 400
rect 78512 0 78568 400
rect 79408 0 79464 400
rect 80304 0 80360 400
rect 81200 0 81256 400
rect 82096 0 82152 400
rect 82992 0 83048 400
rect 83888 0 83944 400
rect 84784 0 84840 400
rect 85680 0 85736 400
rect 86576 0 86632 400
rect 87472 0 87528 400
rect 88368 0 88424 400
rect 89264 0 89320 400
rect 90160 0 90216 400
rect 91056 0 91112 400
rect 91952 0 92008 400
rect 92848 0 92904 400
rect 93744 0 93800 400
rect 94640 0 94696 400
rect 95536 0 95592 400
rect 96432 0 96488 400
rect 97328 0 97384 400
rect 98224 0 98280 400
rect 99120 0 99176 400
rect 100016 0 100072 400
rect 100912 0 100968 400
rect 101808 0 101864 400
rect 102704 0 102760 400
rect 103600 0 103656 400
rect 104496 0 104552 400
rect 105392 0 105448 400
rect 106288 0 106344 400
rect 107184 0 107240 400
rect 108080 0 108136 400
rect 108976 0 109032 400
rect 109872 0 109928 400
rect 110768 0 110824 400
rect 111664 0 111720 400
rect 112560 0 112616 400
rect 113456 0 113512 400
rect 114352 0 114408 400
rect 115248 0 115304 400
rect 116144 0 116200 400
rect 117040 0 117096 400
rect 117936 0 117992 400
rect 118832 0 118888 400
rect 119728 0 119784 400
rect 120624 0 120680 400
rect 121520 0 121576 400
rect 122416 0 122472 400
rect 123312 0 123368 400
rect 124208 0 124264 400
rect 125104 0 125160 400
rect 126000 0 126056 400
rect 126896 0 126952 400
rect 127792 0 127848 400
rect 128688 0 128744 400
rect 129584 0 129640 400
rect 130480 0 130536 400
rect 131376 0 131432 400
rect 132272 0 132328 400
rect 133168 0 133224 400
rect 134064 0 134120 400
rect 134960 0 135016 400
rect 135856 0 135912 400
rect 136752 0 136808 400
rect 137648 0 137704 400
rect 138544 0 138600 400
rect 139440 0 139496 400
rect 140336 0 140392 400
rect 141232 0 141288 400
rect 142128 0 142184 400
rect 143024 0 143080 400
rect 143920 0 143976 400
rect 144816 0 144872 400
rect 145712 0 145768 400
rect 146608 0 146664 400
rect 147504 0 147560 400
rect 148400 0 148456 400
rect 149296 0 149352 400
rect 150192 0 150248 400
rect 151088 0 151144 400
rect 151984 0 152040 400
rect 152880 0 152936 400
rect 153776 0 153832 400
rect 154672 0 154728 400
rect 155568 0 155624 400
rect 156464 0 156520 400
rect 157360 0 157416 400
rect 158256 0 158312 400
rect 159152 0 159208 400
rect 160048 0 160104 400
rect 160944 0 161000 400
rect 161840 0 161896 400
rect 162736 0 162792 400
rect 163632 0 163688 400
rect 164528 0 164584 400
rect 165424 0 165480 400
rect 166320 0 166376 400
rect 167216 0 167272 400
rect 168112 0 168168 400
rect 169008 0 169064 400
rect 169904 0 169960 400
rect 170800 0 170856 400
rect 171696 0 171752 400
rect 172592 0 172648 400
rect 173488 0 173544 400
rect 174384 0 174440 400
rect 175280 0 175336 400
rect 176176 0 176232 400
rect 177072 0 177128 400
rect 177968 0 178024 400
rect 178864 0 178920 400
rect 179760 0 179816 400
rect 180656 0 180712 400
rect 181552 0 181608 400
rect 182448 0 182504 400
rect 183344 0 183400 400
rect 184240 0 184296 400
rect 185136 0 185192 400
rect 186032 0 186088 400
rect 186928 0 186984 400
rect 187824 0 187880 400
rect 188720 0 188776 400
rect 189616 0 189672 400
rect 190512 0 190568 400
rect 191408 0 191464 400
rect 192304 0 192360 400
rect 193200 0 193256 400
rect 194096 0 194152 400
rect 194992 0 195048 400
rect 195888 0 195944 400
rect 196784 0 196840 400
rect 197680 0 197736 400
rect 198576 0 198632 400
rect 199472 0 199528 400
rect 200368 0 200424 400
rect 201264 0 201320 400
rect 202160 0 202216 400
rect 203056 0 203112 400
rect 203952 0 204008 400
rect 204848 0 204904 400
rect 205744 0 205800 400
rect 206640 0 206696 400
rect 207536 0 207592 400
rect 208432 0 208488 400
rect 209328 0 209384 400
rect 210224 0 210280 400
rect 211120 0 211176 400
rect 212016 0 212072 400
rect 212912 0 212968 400
rect 213808 0 213864 400
rect 214704 0 214760 400
rect 215600 0 215656 400
rect 216496 0 216552 400
rect 217392 0 217448 400
rect 218288 0 218344 400
rect 219184 0 219240 400
rect 220080 0 220136 400
rect 220976 0 221032 400
rect 221872 0 221928 400
rect 222768 0 222824 400
rect 223664 0 223720 400
rect 224560 0 224616 400
rect 225456 0 225512 400
rect 226352 0 226408 400
rect 227248 0 227304 400
rect 228144 0 228200 400
rect 229040 0 229096 400
rect 229936 0 229992 400
rect 230832 0 230888 400
rect 231728 0 231784 400
rect 232624 0 232680 400
rect 233520 0 233576 400
rect 234416 0 234472 400
rect 235312 0 235368 400
rect 236208 0 236264 400
rect 237104 0 237160 400
rect 238000 0 238056 400
rect 238896 0 238952 400
rect 239792 0 239848 400
rect 240688 0 240744 400
rect 241584 0 241640 400
rect 242480 0 242536 400
rect 243376 0 243432 400
rect 244272 0 244328 400
rect 245168 0 245224 400
rect 246064 0 246120 400
rect 246960 0 247016 400
rect 247856 0 247912 400
rect 248752 0 248808 400
rect 249648 0 249704 400
rect 250544 0 250600 400
rect 251440 0 251496 400
rect 252336 0 252392 400
rect 253232 0 253288 400
rect 254128 0 254184 400
rect 255024 0 255080 400
rect 255920 0 255976 400
rect 256816 0 256872 400
rect 257712 0 257768 400
rect 258608 0 258664 400
rect 259504 0 259560 400
rect 260400 0 260456 400
rect 261296 0 261352 400
rect 262192 0 262248 400
rect 263088 0 263144 400
rect 263984 0 264040 400
rect 264880 0 264936 400
rect 265776 0 265832 400
rect 266672 0 266728 400
rect 267568 0 267624 400
rect 268464 0 268520 400
rect 269360 0 269416 400
rect 270256 0 270312 400
rect 271152 0 271208 400
rect 272048 0 272104 400
rect 272944 0 273000 400
rect 273840 0 273896 400
rect 274736 0 274792 400
rect 275632 0 275688 400
rect 276528 0 276584 400
rect 277424 0 277480 400
rect 278320 0 278376 400
<< obsm2 >>
rect 462 288409 4226 288439
rect 4342 288409 12178 288439
rect 12294 288409 20130 288439
rect 20246 288409 28082 288439
rect 28198 288409 36034 288439
rect 36150 288409 43986 288439
rect 44102 288409 51938 288439
rect 52054 288409 59890 288439
rect 60006 288409 67842 288439
rect 67958 288409 75794 288439
rect 75910 288409 83746 288439
rect 83862 288409 91698 288439
rect 91814 288409 99650 288439
rect 99766 288409 107602 288439
rect 107718 288409 115554 288439
rect 115670 288409 123506 288439
rect 123622 288409 131458 288439
rect 131574 288409 139410 288439
rect 139526 288409 147362 288439
rect 147478 288409 155314 288439
rect 155430 288409 163266 288439
rect 163382 288409 171218 288439
rect 171334 288409 179170 288439
rect 179286 288409 187122 288439
rect 187238 288409 195074 288439
rect 195190 288409 203026 288439
rect 203142 288409 210978 288439
rect 211094 288409 218930 288439
rect 219046 288409 226882 288439
rect 226998 288409 234834 288439
rect 234950 288409 242786 288439
rect 242902 288409 250738 288439
rect 250854 288409 258690 288439
rect 258806 288409 266642 288439
rect 266758 288409 274594 288439
rect 274710 288409 282546 288439
rect 282662 288409 286370 288439
rect 462 430 286370 288409
rect 462 289 8594 430
rect 8710 289 9490 430
rect 9606 289 10386 430
rect 10502 289 11282 430
rect 11398 289 12178 430
rect 12294 289 13074 430
rect 13190 289 13970 430
rect 14086 289 14866 430
rect 14982 289 15762 430
rect 15878 289 16658 430
rect 16774 289 17554 430
rect 17670 289 18450 430
rect 18566 289 19346 430
rect 19462 289 20242 430
rect 20358 289 21138 430
rect 21254 289 22034 430
rect 22150 289 22930 430
rect 23046 289 23826 430
rect 23942 289 24722 430
rect 24838 289 25618 430
rect 25734 289 26514 430
rect 26630 289 27410 430
rect 27526 289 28306 430
rect 28422 289 29202 430
rect 29318 289 30098 430
rect 30214 289 30994 430
rect 31110 289 31890 430
rect 32006 289 32786 430
rect 32902 289 33682 430
rect 33798 289 34578 430
rect 34694 289 35474 430
rect 35590 289 36370 430
rect 36486 289 37266 430
rect 37382 289 38162 430
rect 38278 289 39058 430
rect 39174 289 39954 430
rect 40070 289 40850 430
rect 40966 289 41746 430
rect 41862 289 42642 430
rect 42758 289 43538 430
rect 43654 289 44434 430
rect 44550 289 45330 430
rect 45446 289 46226 430
rect 46342 289 47122 430
rect 47238 289 48018 430
rect 48134 289 48914 430
rect 49030 289 49810 430
rect 49926 289 50706 430
rect 50822 289 51602 430
rect 51718 289 52498 430
rect 52614 289 53394 430
rect 53510 289 54290 430
rect 54406 289 55186 430
rect 55302 289 56082 430
rect 56198 289 56978 430
rect 57094 289 57874 430
rect 57990 289 58770 430
rect 58886 289 59666 430
rect 59782 289 60562 430
rect 60678 289 61458 430
rect 61574 289 62354 430
rect 62470 289 63250 430
rect 63366 289 64146 430
rect 64262 289 65042 430
rect 65158 289 65938 430
rect 66054 289 66834 430
rect 66950 289 67730 430
rect 67846 289 68626 430
rect 68742 289 69522 430
rect 69638 289 70418 430
rect 70534 289 71314 430
rect 71430 289 72210 430
rect 72326 289 73106 430
rect 73222 289 74002 430
rect 74118 289 74898 430
rect 75014 289 75794 430
rect 75910 289 76690 430
rect 76806 289 77586 430
rect 77702 289 78482 430
rect 78598 289 79378 430
rect 79494 289 80274 430
rect 80390 289 81170 430
rect 81286 289 82066 430
rect 82182 289 82962 430
rect 83078 289 83858 430
rect 83974 289 84754 430
rect 84870 289 85650 430
rect 85766 289 86546 430
rect 86662 289 87442 430
rect 87558 289 88338 430
rect 88454 289 89234 430
rect 89350 289 90130 430
rect 90246 289 91026 430
rect 91142 289 91922 430
rect 92038 289 92818 430
rect 92934 289 93714 430
rect 93830 289 94610 430
rect 94726 289 95506 430
rect 95622 289 96402 430
rect 96518 289 97298 430
rect 97414 289 98194 430
rect 98310 289 99090 430
rect 99206 289 99986 430
rect 100102 289 100882 430
rect 100998 289 101778 430
rect 101894 289 102674 430
rect 102790 289 103570 430
rect 103686 289 104466 430
rect 104582 289 105362 430
rect 105478 289 106258 430
rect 106374 289 107154 430
rect 107270 289 108050 430
rect 108166 289 108946 430
rect 109062 289 109842 430
rect 109958 289 110738 430
rect 110854 289 111634 430
rect 111750 289 112530 430
rect 112646 289 113426 430
rect 113542 289 114322 430
rect 114438 289 115218 430
rect 115334 289 116114 430
rect 116230 289 117010 430
rect 117126 289 117906 430
rect 118022 289 118802 430
rect 118918 289 119698 430
rect 119814 289 120594 430
rect 120710 289 121490 430
rect 121606 289 122386 430
rect 122502 289 123282 430
rect 123398 289 124178 430
rect 124294 289 125074 430
rect 125190 289 125970 430
rect 126086 289 126866 430
rect 126982 289 127762 430
rect 127878 289 128658 430
rect 128774 289 129554 430
rect 129670 289 130450 430
rect 130566 289 131346 430
rect 131462 289 132242 430
rect 132358 289 133138 430
rect 133254 289 134034 430
rect 134150 289 134930 430
rect 135046 289 135826 430
rect 135942 289 136722 430
rect 136838 289 137618 430
rect 137734 289 138514 430
rect 138630 289 139410 430
rect 139526 289 140306 430
rect 140422 289 141202 430
rect 141318 289 142098 430
rect 142214 289 142994 430
rect 143110 289 143890 430
rect 144006 289 144786 430
rect 144902 289 145682 430
rect 145798 289 146578 430
rect 146694 289 147474 430
rect 147590 289 148370 430
rect 148486 289 149266 430
rect 149382 289 150162 430
rect 150278 289 151058 430
rect 151174 289 151954 430
rect 152070 289 152850 430
rect 152966 289 153746 430
rect 153862 289 154642 430
rect 154758 289 155538 430
rect 155654 289 156434 430
rect 156550 289 157330 430
rect 157446 289 158226 430
rect 158342 289 159122 430
rect 159238 289 160018 430
rect 160134 289 160914 430
rect 161030 289 161810 430
rect 161926 289 162706 430
rect 162822 289 163602 430
rect 163718 289 164498 430
rect 164614 289 165394 430
rect 165510 289 166290 430
rect 166406 289 167186 430
rect 167302 289 168082 430
rect 168198 289 168978 430
rect 169094 289 169874 430
rect 169990 289 170770 430
rect 170886 289 171666 430
rect 171782 289 172562 430
rect 172678 289 173458 430
rect 173574 289 174354 430
rect 174470 289 175250 430
rect 175366 289 176146 430
rect 176262 289 177042 430
rect 177158 289 177938 430
rect 178054 289 178834 430
rect 178950 289 179730 430
rect 179846 289 180626 430
rect 180742 289 181522 430
rect 181638 289 182418 430
rect 182534 289 183314 430
rect 183430 289 184210 430
rect 184326 289 185106 430
rect 185222 289 186002 430
rect 186118 289 186898 430
rect 187014 289 187794 430
rect 187910 289 188690 430
rect 188806 289 189586 430
rect 189702 289 190482 430
rect 190598 289 191378 430
rect 191494 289 192274 430
rect 192390 289 193170 430
rect 193286 289 194066 430
rect 194182 289 194962 430
rect 195078 289 195858 430
rect 195974 289 196754 430
rect 196870 289 197650 430
rect 197766 289 198546 430
rect 198662 289 199442 430
rect 199558 289 200338 430
rect 200454 289 201234 430
rect 201350 289 202130 430
rect 202246 289 203026 430
rect 203142 289 203922 430
rect 204038 289 204818 430
rect 204934 289 205714 430
rect 205830 289 206610 430
rect 206726 289 207506 430
rect 207622 289 208402 430
rect 208518 289 209298 430
rect 209414 289 210194 430
rect 210310 289 211090 430
rect 211206 289 211986 430
rect 212102 289 212882 430
rect 212998 289 213778 430
rect 213894 289 214674 430
rect 214790 289 215570 430
rect 215686 289 216466 430
rect 216582 289 217362 430
rect 217478 289 218258 430
rect 218374 289 219154 430
rect 219270 289 220050 430
rect 220166 289 220946 430
rect 221062 289 221842 430
rect 221958 289 222738 430
rect 222854 289 223634 430
rect 223750 289 224530 430
rect 224646 289 225426 430
rect 225542 289 226322 430
rect 226438 289 227218 430
rect 227334 289 228114 430
rect 228230 289 229010 430
rect 229126 289 229906 430
rect 230022 289 230802 430
rect 230918 289 231698 430
rect 231814 289 232594 430
rect 232710 289 233490 430
rect 233606 289 234386 430
rect 234502 289 235282 430
rect 235398 289 236178 430
rect 236294 289 237074 430
rect 237190 289 237970 430
rect 238086 289 238866 430
rect 238982 289 239762 430
rect 239878 289 240658 430
rect 240774 289 241554 430
rect 241670 289 242450 430
rect 242566 289 243346 430
rect 243462 289 244242 430
rect 244358 289 245138 430
rect 245254 289 246034 430
rect 246150 289 246930 430
rect 247046 289 247826 430
rect 247942 289 248722 430
rect 248838 289 249618 430
rect 249734 289 250514 430
rect 250630 289 251410 430
rect 251526 289 252306 430
rect 252422 289 253202 430
rect 253318 289 254098 430
rect 254214 289 254994 430
rect 255110 289 255890 430
rect 256006 289 256786 430
rect 256902 289 257682 430
rect 257798 289 258578 430
rect 258694 289 259474 430
rect 259590 289 260370 430
rect 260486 289 261266 430
rect 261382 289 262162 430
rect 262278 289 263058 430
rect 263174 289 263954 430
rect 264070 289 264850 430
rect 264966 289 265746 430
rect 265862 289 266642 430
rect 266758 289 267538 430
rect 267654 289 268434 430
rect 268550 289 269330 430
rect 269446 289 270226 430
rect 270342 289 271122 430
rect 271238 289 272018 430
rect 272134 289 272914 430
rect 273030 289 273810 430
rect 273926 289 274706 430
rect 274822 289 275602 430
rect 275718 289 276498 430
rect 276614 289 277394 430
rect 277510 289 278290 430
rect 278406 289 286370 430
<< metal3 >>
rect 286647 284144 287047 284200
rect 0 283808 400 283864
rect 286647 278768 287047 278824
rect 0 278544 400 278600
rect 286647 273392 287047 273448
rect 0 273280 400 273336
rect 0 268016 400 268072
rect 286647 268016 287047 268072
rect 0 262752 400 262808
rect 286647 262640 287047 262696
rect 0 257488 400 257544
rect 286647 257264 287047 257320
rect 0 252224 400 252280
rect 286647 251888 287047 251944
rect 0 246960 400 247016
rect 286647 246512 287047 246568
rect 0 241696 400 241752
rect 286647 241136 287047 241192
rect 0 236432 400 236488
rect 286647 235760 287047 235816
rect 0 231168 400 231224
rect 286647 230384 287047 230440
rect 0 225904 400 225960
rect 286647 225008 287047 225064
rect 0 220640 400 220696
rect 286647 219632 287047 219688
rect 0 215376 400 215432
rect 286647 214256 287047 214312
rect 0 210112 400 210168
rect 286647 208880 287047 208936
rect 0 204848 400 204904
rect 286647 203504 287047 203560
rect 0 199584 400 199640
rect 286647 198128 287047 198184
rect 0 194320 400 194376
rect 286647 192752 287047 192808
rect 0 189056 400 189112
rect 286647 187376 287047 187432
rect 0 183792 400 183848
rect 286647 182000 287047 182056
rect 0 178528 400 178584
rect 286647 176624 287047 176680
rect 0 173264 400 173320
rect 286647 171248 287047 171304
rect 0 168000 400 168056
rect 286647 165872 287047 165928
rect 0 162736 400 162792
rect 286647 160496 287047 160552
rect 0 157472 400 157528
rect 286647 155120 287047 155176
rect 0 152208 400 152264
rect 286647 149744 287047 149800
rect 0 146944 400 147000
rect 286647 144368 287047 144424
rect 0 141680 400 141736
rect 286647 138992 287047 139048
rect 0 136416 400 136472
rect 286647 133616 287047 133672
rect 0 131152 400 131208
rect 286647 128240 287047 128296
rect 0 125888 400 125944
rect 286647 122864 287047 122920
rect 0 120624 400 120680
rect 286647 117488 287047 117544
rect 0 115360 400 115416
rect 286647 112112 287047 112168
rect 0 110096 400 110152
rect 286647 106736 287047 106792
rect 0 104832 400 104888
rect 286647 101360 287047 101416
rect 0 99568 400 99624
rect 286647 95984 287047 96040
rect 0 94304 400 94360
rect 286647 90608 287047 90664
rect 0 89040 400 89096
rect 286647 85232 287047 85288
rect 0 83776 400 83832
rect 286647 79856 287047 79912
rect 0 78512 400 78568
rect 286647 74480 287047 74536
rect 0 73248 400 73304
rect 286647 69104 287047 69160
rect 0 67984 400 68040
rect 286647 63728 287047 63784
rect 0 62720 400 62776
rect 286647 58352 287047 58408
rect 0 57456 400 57512
rect 286647 52976 287047 53032
rect 0 52192 400 52248
rect 286647 47600 287047 47656
rect 0 46928 400 46984
rect 286647 42224 287047 42280
rect 0 41664 400 41720
rect 286647 36848 287047 36904
rect 0 36400 400 36456
rect 286647 31472 287047 31528
rect 0 31136 400 31192
rect 286647 26096 287047 26152
rect 0 25872 400 25928
rect 286647 20720 287047 20776
rect 0 20608 400 20664
rect 0 15344 400 15400
rect 286647 15344 287047 15400
rect 0 10080 400 10136
rect 286647 9968 287047 10024
rect 0 4816 400 4872
rect 286647 4592 287047 4648
<< obsm3 >>
rect 400 284230 286647 287434
rect 400 284114 286617 284230
rect 400 283894 286647 284114
rect 430 283778 286647 283894
rect 400 278854 286647 283778
rect 400 278738 286617 278854
rect 400 278630 286647 278738
rect 430 278514 286647 278630
rect 400 273478 286647 278514
rect 400 273366 286617 273478
rect 430 273362 286617 273366
rect 430 273250 286647 273362
rect 400 268102 286647 273250
rect 430 267986 286617 268102
rect 400 262838 286647 267986
rect 430 262726 286647 262838
rect 430 262722 286617 262726
rect 400 262610 286617 262722
rect 400 257574 286647 262610
rect 430 257458 286647 257574
rect 400 257350 286647 257458
rect 400 257234 286617 257350
rect 400 252310 286647 257234
rect 430 252194 286647 252310
rect 400 251974 286647 252194
rect 400 251858 286617 251974
rect 400 247046 286647 251858
rect 430 246930 286647 247046
rect 400 246598 286647 246930
rect 400 246482 286617 246598
rect 400 241782 286647 246482
rect 430 241666 286647 241782
rect 400 241222 286647 241666
rect 400 241106 286617 241222
rect 400 236518 286647 241106
rect 430 236402 286647 236518
rect 400 235846 286647 236402
rect 400 235730 286617 235846
rect 400 231254 286647 235730
rect 430 231138 286647 231254
rect 400 230470 286647 231138
rect 400 230354 286617 230470
rect 400 225990 286647 230354
rect 430 225874 286647 225990
rect 400 225094 286647 225874
rect 400 224978 286617 225094
rect 400 220726 286647 224978
rect 430 220610 286647 220726
rect 400 219718 286647 220610
rect 400 219602 286617 219718
rect 400 215462 286647 219602
rect 430 215346 286647 215462
rect 400 214342 286647 215346
rect 400 214226 286617 214342
rect 400 210198 286647 214226
rect 430 210082 286647 210198
rect 400 208966 286647 210082
rect 400 208850 286617 208966
rect 400 204934 286647 208850
rect 430 204818 286647 204934
rect 400 203590 286647 204818
rect 400 203474 286617 203590
rect 400 199670 286647 203474
rect 430 199554 286647 199670
rect 400 198214 286647 199554
rect 400 198098 286617 198214
rect 400 194406 286647 198098
rect 430 194290 286647 194406
rect 400 192838 286647 194290
rect 400 192722 286617 192838
rect 400 189142 286647 192722
rect 430 189026 286647 189142
rect 400 187462 286647 189026
rect 400 187346 286617 187462
rect 400 183878 286647 187346
rect 430 183762 286647 183878
rect 400 182086 286647 183762
rect 400 181970 286617 182086
rect 400 178614 286647 181970
rect 430 178498 286647 178614
rect 400 176710 286647 178498
rect 400 176594 286617 176710
rect 400 173350 286647 176594
rect 430 173234 286647 173350
rect 400 171334 286647 173234
rect 400 171218 286617 171334
rect 400 168086 286647 171218
rect 430 167970 286647 168086
rect 400 165958 286647 167970
rect 400 165842 286617 165958
rect 400 162822 286647 165842
rect 430 162706 286647 162822
rect 400 160582 286647 162706
rect 400 160466 286617 160582
rect 400 157558 286647 160466
rect 430 157442 286647 157558
rect 400 155206 286647 157442
rect 400 155090 286617 155206
rect 400 152294 286647 155090
rect 430 152178 286647 152294
rect 400 149830 286647 152178
rect 400 149714 286617 149830
rect 400 147030 286647 149714
rect 430 146914 286647 147030
rect 400 144454 286647 146914
rect 400 144338 286617 144454
rect 400 141766 286647 144338
rect 430 141650 286647 141766
rect 400 139078 286647 141650
rect 400 138962 286617 139078
rect 400 136502 286647 138962
rect 430 136386 286647 136502
rect 400 133702 286647 136386
rect 400 133586 286617 133702
rect 400 131238 286647 133586
rect 430 131122 286647 131238
rect 400 128326 286647 131122
rect 400 128210 286617 128326
rect 400 125974 286647 128210
rect 430 125858 286647 125974
rect 400 122950 286647 125858
rect 400 122834 286617 122950
rect 400 120710 286647 122834
rect 430 120594 286647 120710
rect 400 117574 286647 120594
rect 400 117458 286617 117574
rect 400 115446 286647 117458
rect 430 115330 286647 115446
rect 400 112198 286647 115330
rect 400 112082 286617 112198
rect 400 110182 286647 112082
rect 430 110066 286647 110182
rect 400 106822 286647 110066
rect 400 106706 286617 106822
rect 400 104918 286647 106706
rect 430 104802 286647 104918
rect 400 101446 286647 104802
rect 400 101330 286617 101446
rect 400 99654 286647 101330
rect 430 99538 286647 99654
rect 400 96070 286647 99538
rect 400 95954 286617 96070
rect 400 94390 286647 95954
rect 430 94274 286647 94390
rect 400 90694 286647 94274
rect 400 90578 286617 90694
rect 400 89126 286647 90578
rect 430 89010 286647 89126
rect 400 85318 286647 89010
rect 400 85202 286617 85318
rect 400 83862 286647 85202
rect 430 83746 286647 83862
rect 400 79942 286647 83746
rect 400 79826 286617 79942
rect 400 78598 286647 79826
rect 430 78482 286647 78598
rect 400 74566 286647 78482
rect 400 74450 286617 74566
rect 400 73334 286647 74450
rect 430 73218 286647 73334
rect 400 69190 286647 73218
rect 400 69074 286617 69190
rect 400 68070 286647 69074
rect 430 67954 286647 68070
rect 400 63814 286647 67954
rect 400 63698 286617 63814
rect 400 62806 286647 63698
rect 430 62690 286647 62806
rect 400 58438 286647 62690
rect 400 58322 286617 58438
rect 400 57542 286647 58322
rect 430 57426 286647 57542
rect 400 53062 286647 57426
rect 400 52946 286617 53062
rect 400 52278 286647 52946
rect 430 52162 286647 52278
rect 400 47686 286647 52162
rect 400 47570 286617 47686
rect 400 47014 286647 47570
rect 430 46898 286647 47014
rect 400 42310 286647 46898
rect 400 42194 286617 42310
rect 400 41750 286647 42194
rect 430 41634 286647 41750
rect 400 36934 286647 41634
rect 400 36818 286617 36934
rect 400 36486 286647 36818
rect 430 36370 286647 36486
rect 400 31558 286647 36370
rect 400 31442 286617 31558
rect 400 31222 286647 31442
rect 430 31106 286647 31222
rect 400 26182 286647 31106
rect 400 26066 286617 26182
rect 400 25958 286647 26066
rect 430 25842 286647 25958
rect 400 20806 286647 25842
rect 400 20694 286617 20806
rect 430 20690 286617 20694
rect 430 20578 286647 20690
rect 400 15430 286647 20578
rect 430 15314 286617 15430
rect 400 10166 286647 15314
rect 430 10054 286647 10166
rect 430 10050 286617 10054
rect 400 9938 286617 10050
rect 400 4902 286647 9938
rect 430 4786 286647 4902
rect 400 4678 286647 4786
rect 400 4562 286617 4678
rect 400 294 286647 4562
<< metal4 >>
rect 2224 1538 2384 286974
rect 9904 1538 10064 286974
rect 17584 1538 17744 286974
rect 25264 1538 25424 286974
rect 32944 1538 33104 286974
rect 40624 1538 40784 286974
rect 48304 1538 48464 286974
rect 55984 1538 56144 286974
rect 63664 1538 63824 286974
rect 71344 1538 71504 286974
rect 79024 1538 79184 286974
rect 86704 1538 86864 286974
rect 94384 1538 94544 286974
rect 102064 1538 102224 286974
rect 109744 1538 109904 286974
rect 117424 1538 117584 286974
rect 125104 1538 125264 286974
rect 132784 1538 132944 286974
rect 140464 1538 140624 286974
rect 148144 1538 148304 286974
rect 155824 1538 155984 286974
rect 163504 1538 163664 286974
rect 171184 1538 171344 286974
rect 178864 1538 179024 286974
rect 186544 1538 186704 286974
rect 194224 1538 194384 286974
rect 201904 1538 202064 286974
rect 209584 1538 209744 286974
rect 217264 1538 217424 286974
rect 224944 1538 225104 286974
rect 232624 1538 232784 286974
rect 240304 1538 240464 286974
rect 247984 1538 248144 286974
rect 255664 1538 255824 286974
rect 263344 1538 263504 286974
rect 271024 1538 271184 286974
rect 278704 1538 278864 286974
<< obsm4 >>
rect 1022 287004 285586 287439
rect 1022 1508 2194 287004
rect 2414 1508 9874 287004
rect 10094 1508 17554 287004
rect 17774 1508 25234 287004
rect 25454 1508 32914 287004
rect 33134 1508 40594 287004
rect 40814 1508 48274 287004
rect 48494 1508 55954 287004
rect 56174 1508 63634 287004
rect 63854 1508 71314 287004
rect 71534 1508 78994 287004
rect 79214 1508 86674 287004
rect 86894 1508 94354 287004
rect 94574 1508 102034 287004
rect 102254 1508 109714 287004
rect 109934 1508 117394 287004
rect 117614 1508 125074 287004
rect 125294 1508 132754 287004
rect 132974 1508 140434 287004
rect 140654 1508 148114 287004
rect 148334 1508 155794 287004
rect 156014 1508 163474 287004
rect 163694 1508 171154 287004
rect 171374 1508 178834 287004
rect 179054 1508 186514 287004
rect 186734 1508 194194 287004
rect 194414 1508 201874 287004
rect 202094 1508 209554 287004
rect 209774 1508 217234 287004
rect 217454 1508 224914 287004
rect 225134 1508 232594 287004
rect 232814 1508 240274 287004
rect 240494 1508 247954 287004
rect 248174 1508 255634 287004
rect 255854 1508 263314 287004
rect 263534 1508 270994 287004
rect 271214 1508 278674 287004
rect 278894 1508 285586 287004
rect 1022 681 285586 1508
<< labels >>
rlabel metal3 s 286647 117488 287047 117544 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 218960 288439 219016 288839 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 187152 288439 187208 288839 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 155344 288439 155400 288839 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 123536 288439 123592 288839 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 91728 288439 91784 288839 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 59920 288439 59976 288839 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 28112 288439 28168 288839 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s 0 283808 400 283864 6 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s 0 262752 400 262808 6 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s 0 241696 400 241752 6 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 286647 138992 287047 139048 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s 0 220640 400 220696 6 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s 0 199584 400 199640 6 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s 0 178528 400 178584 6 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s 0 157472 400 157528 6 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s 0 136416 400 136472 6 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s 0 115360 400 115416 6 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s 0 94304 400 94360 6 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s 0 73248 400 73304 6 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s 0 52192 400 52248 6 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 286647 160496 287047 160552 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 286647 182000 287047 182056 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 286647 203504 287047 203560 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 286647 225008 287047 225064 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 286647 246512 287047 246568 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 286647 268016 287047 268072 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 282576 288439 282632 288839 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 250768 288439 250824 288839 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 286647 4592 287047 4648 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 286647 187376 287047 187432 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 286647 208880 287047 208936 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 286647 230384 287047 230440 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 286647 251888 287047 251944 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 286647 273392 287047 273448 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 274624 288439 274680 288839 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 242816 288439 242872 288839 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 211008 288439 211064 288839 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 179200 288439 179256 288839 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 147392 288439 147448 288839 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 286647 20720 287047 20776 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 115584 288439 115640 288839 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 83776 288439 83832 288839 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 51968 288439 52024 288839 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 20160 288439 20216 288839 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s 0 278544 400 278600 6 io_in[24]
port 46 nsew signal input
rlabel metal3 s 0 257488 400 257544 6 io_in[25]
port 47 nsew signal input
rlabel metal3 s 0 236432 400 236488 6 io_in[26]
port 48 nsew signal input
rlabel metal3 s 0 215376 400 215432 6 io_in[27]
port 49 nsew signal input
rlabel metal3 s 0 194320 400 194376 6 io_in[28]
port 50 nsew signal input
rlabel metal3 s 0 173264 400 173320 6 io_in[29]
port 51 nsew signal input
rlabel metal3 s 286647 36848 287047 36904 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s 0 152208 400 152264 6 io_in[30]
port 53 nsew signal input
rlabel metal3 s 0 131152 400 131208 6 io_in[31]
port 54 nsew signal input
rlabel metal3 s 0 110096 400 110152 6 io_in[32]
port 55 nsew signal input
rlabel metal3 s 0 89040 400 89096 6 io_in[33]
port 56 nsew signal input
rlabel metal3 s 0 67984 400 68040 6 io_in[34]
port 57 nsew signal input
rlabel metal3 s 0 46928 400 46984 6 io_in[35]
port 58 nsew signal input
rlabel metal3 s 0 31136 400 31192 6 io_in[36]
port 59 nsew signal input
rlabel metal3 s 0 15344 400 15400 6 io_in[37]
port 60 nsew signal input
rlabel metal3 s 286647 52976 287047 53032 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 286647 69104 287047 69160 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 286647 85232 287047 85288 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 286647 101360 287047 101416 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 286647 122864 287047 122920 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 286647 144368 287047 144424 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 286647 165872 287047 165928 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 286647 15344 287047 15400 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 286647 198128 287047 198184 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 286647 219632 287047 219688 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 286647 241136 287047 241192 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 286647 262640 287047 262696 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 286647 284144 287047 284200 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 258720 288439 258776 288839 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 226912 288439 226968 288839 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 195104 288439 195160 288839 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 163296 288439 163352 288839 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 131488 288439 131544 288839 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 286647 31472 287047 31528 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 99680 288439 99736 288839 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 67872 288439 67928 288839 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 36064 288439 36120 288839 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 4256 288439 4312 288839 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s 0 268016 400 268072 6 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s 0 246960 400 247016 6 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s 0 225904 400 225960 6 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s 0 204848 400 204904 6 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s 0 183792 400 183848 6 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s 0 162736 400 162792 6 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 286647 47600 287047 47656 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s 0 141680 400 141736 6 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s 0 120624 400 120680 6 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s 0 99568 400 99624 6 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s 0 78512 400 78568 6 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s 0 57456 400 57512 6 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s 0 36400 400 36456 6 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s 0 20608 400 20664 6 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s 0 4816 400 4872 6 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 286647 63728 287047 63784 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 286647 79856 287047 79912 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 286647 95984 287047 96040 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 286647 112112 287047 112168 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 286647 133616 287047 133672 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 286647 155120 287047 155176 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 286647 176624 287047 176680 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 286647 9968 287047 10024 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 286647 192752 287047 192808 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 286647 214256 287047 214312 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 286647 235760 287047 235816 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 286647 257264 287047 257320 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 286647 278768 287047 278824 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 266672 288439 266728 288839 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 234864 288439 234920 288839 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 203056 288439 203112 288839 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 171248 288439 171304 288839 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 139440 288439 139496 288839 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 286647 26096 287047 26152 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 107632 288439 107688 288839 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 75824 288439 75880 288839 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 44016 288439 44072 288839 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 12208 288439 12264 288839 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s 0 273280 400 273336 6 io_out[24]
port 122 nsew signal output
rlabel metal3 s 0 252224 400 252280 6 io_out[25]
port 123 nsew signal output
rlabel metal3 s 0 231168 400 231224 6 io_out[26]
port 124 nsew signal output
rlabel metal3 s 0 210112 400 210168 6 io_out[27]
port 125 nsew signal output
rlabel metal3 s 0 189056 400 189112 6 io_out[28]
port 126 nsew signal output
rlabel metal3 s 0 168000 400 168056 6 io_out[29]
port 127 nsew signal output
rlabel metal3 s 286647 42224 287047 42280 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s 0 146944 400 147000 6 io_out[30]
port 129 nsew signal output
rlabel metal3 s 0 125888 400 125944 6 io_out[31]
port 130 nsew signal output
rlabel metal3 s 0 104832 400 104888 6 io_out[32]
port 131 nsew signal output
rlabel metal3 s 0 83776 400 83832 6 io_out[33]
port 132 nsew signal output
rlabel metal3 s 0 62720 400 62776 6 io_out[34]
port 133 nsew signal output
rlabel metal3 s 0 41664 400 41720 6 io_out[35]
port 134 nsew signal output
rlabel metal3 s 0 25872 400 25928 6 io_out[36]
port 135 nsew signal output
rlabel metal3 s 0 10080 400 10136 6 io_out[37]
port 136 nsew signal output
rlabel metal3 s 286647 58352 287047 58408 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 286647 74480 287047 74536 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 286647 90608 287047 90664 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 286647 106736 287047 106792 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 286647 128240 287047 128296 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 286647 149744 287047 149800 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 286647 171248 287047 171304 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 103600 0 103656 400 6 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 130480 0 130536 400 6 la_data_in[10]
port 145 nsew signal input
rlabel metal2 s 133168 0 133224 400 6 la_data_in[11]
port 146 nsew signal input
rlabel metal2 s 135856 0 135912 400 6 la_data_in[12]
port 147 nsew signal input
rlabel metal2 s 138544 0 138600 400 6 la_data_in[13]
port 148 nsew signal input
rlabel metal2 s 141232 0 141288 400 6 la_data_in[14]
port 149 nsew signal input
rlabel metal2 s 143920 0 143976 400 6 la_data_in[15]
port 150 nsew signal input
rlabel metal2 s 146608 0 146664 400 6 la_data_in[16]
port 151 nsew signal input
rlabel metal2 s 149296 0 149352 400 6 la_data_in[17]
port 152 nsew signal input
rlabel metal2 s 151984 0 152040 400 6 la_data_in[18]
port 153 nsew signal input
rlabel metal2 s 154672 0 154728 400 6 la_data_in[19]
port 154 nsew signal input
rlabel metal2 s 106288 0 106344 400 6 la_data_in[1]
port 155 nsew signal input
rlabel metal2 s 157360 0 157416 400 6 la_data_in[20]
port 156 nsew signal input
rlabel metal2 s 160048 0 160104 400 6 la_data_in[21]
port 157 nsew signal input
rlabel metal2 s 162736 0 162792 400 6 la_data_in[22]
port 158 nsew signal input
rlabel metal2 s 165424 0 165480 400 6 la_data_in[23]
port 159 nsew signal input
rlabel metal2 s 168112 0 168168 400 6 la_data_in[24]
port 160 nsew signal input
rlabel metal2 s 170800 0 170856 400 6 la_data_in[25]
port 161 nsew signal input
rlabel metal2 s 173488 0 173544 400 6 la_data_in[26]
port 162 nsew signal input
rlabel metal2 s 176176 0 176232 400 6 la_data_in[27]
port 163 nsew signal input
rlabel metal2 s 178864 0 178920 400 6 la_data_in[28]
port 164 nsew signal input
rlabel metal2 s 181552 0 181608 400 6 la_data_in[29]
port 165 nsew signal input
rlabel metal2 s 108976 0 109032 400 6 la_data_in[2]
port 166 nsew signal input
rlabel metal2 s 184240 0 184296 400 6 la_data_in[30]
port 167 nsew signal input
rlabel metal2 s 186928 0 186984 400 6 la_data_in[31]
port 168 nsew signal input
rlabel metal2 s 189616 0 189672 400 6 la_data_in[32]
port 169 nsew signal input
rlabel metal2 s 192304 0 192360 400 6 la_data_in[33]
port 170 nsew signal input
rlabel metal2 s 194992 0 195048 400 6 la_data_in[34]
port 171 nsew signal input
rlabel metal2 s 197680 0 197736 400 6 la_data_in[35]
port 172 nsew signal input
rlabel metal2 s 200368 0 200424 400 6 la_data_in[36]
port 173 nsew signal input
rlabel metal2 s 203056 0 203112 400 6 la_data_in[37]
port 174 nsew signal input
rlabel metal2 s 205744 0 205800 400 6 la_data_in[38]
port 175 nsew signal input
rlabel metal2 s 208432 0 208488 400 6 la_data_in[39]
port 176 nsew signal input
rlabel metal2 s 111664 0 111720 400 6 la_data_in[3]
port 177 nsew signal input
rlabel metal2 s 211120 0 211176 400 6 la_data_in[40]
port 178 nsew signal input
rlabel metal2 s 213808 0 213864 400 6 la_data_in[41]
port 179 nsew signal input
rlabel metal2 s 216496 0 216552 400 6 la_data_in[42]
port 180 nsew signal input
rlabel metal2 s 219184 0 219240 400 6 la_data_in[43]
port 181 nsew signal input
rlabel metal2 s 221872 0 221928 400 6 la_data_in[44]
port 182 nsew signal input
rlabel metal2 s 224560 0 224616 400 6 la_data_in[45]
port 183 nsew signal input
rlabel metal2 s 227248 0 227304 400 6 la_data_in[46]
port 184 nsew signal input
rlabel metal2 s 229936 0 229992 400 6 la_data_in[47]
port 185 nsew signal input
rlabel metal2 s 232624 0 232680 400 6 la_data_in[48]
port 186 nsew signal input
rlabel metal2 s 235312 0 235368 400 6 la_data_in[49]
port 187 nsew signal input
rlabel metal2 s 114352 0 114408 400 6 la_data_in[4]
port 188 nsew signal input
rlabel metal2 s 238000 0 238056 400 6 la_data_in[50]
port 189 nsew signal input
rlabel metal2 s 240688 0 240744 400 6 la_data_in[51]
port 190 nsew signal input
rlabel metal2 s 243376 0 243432 400 6 la_data_in[52]
port 191 nsew signal input
rlabel metal2 s 246064 0 246120 400 6 la_data_in[53]
port 192 nsew signal input
rlabel metal2 s 248752 0 248808 400 6 la_data_in[54]
port 193 nsew signal input
rlabel metal2 s 251440 0 251496 400 6 la_data_in[55]
port 194 nsew signal input
rlabel metal2 s 254128 0 254184 400 6 la_data_in[56]
port 195 nsew signal input
rlabel metal2 s 256816 0 256872 400 6 la_data_in[57]
port 196 nsew signal input
rlabel metal2 s 259504 0 259560 400 6 la_data_in[58]
port 197 nsew signal input
rlabel metal2 s 262192 0 262248 400 6 la_data_in[59]
port 198 nsew signal input
rlabel metal2 s 117040 0 117096 400 6 la_data_in[5]
port 199 nsew signal input
rlabel metal2 s 264880 0 264936 400 6 la_data_in[60]
port 200 nsew signal input
rlabel metal2 s 267568 0 267624 400 6 la_data_in[61]
port 201 nsew signal input
rlabel metal2 s 270256 0 270312 400 6 la_data_in[62]
port 202 nsew signal input
rlabel metal2 s 272944 0 273000 400 6 la_data_in[63]
port 203 nsew signal input
rlabel metal2 s 119728 0 119784 400 6 la_data_in[6]
port 204 nsew signal input
rlabel metal2 s 122416 0 122472 400 6 la_data_in[7]
port 205 nsew signal input
rlabel metal2 s 125104 0 125160 400 6 la_data_in[8]
port 206 nsew signal input
rlabel metal2 s 127792 0 127848 400 6 la_data_in[9]
port 207 nsew signal input
rlabel metal2 s 104496 0 104552 400 6 la_data_out[0]
port 208 nsew signal output
rlabel metal2 s 131376 0 131432 400 6 la_data_out[10]
port 209 nsew signal output
rlabel metal2 s 134064 0 134120 400 6 la_data_out[11]
port 210 nsew signal output
rlabel metal2 s 136752 0 136808 400 6 la_data_out[12]
port 211 nsew signal output
rlabel metal2 s 139440 0 139496 400 6 la_data_out[13]
port 212 nsew signal output
rlabel metal2 s 142128 0 142184 400 6 la_data_out[14]
port 213 nsew signal output
rlabel metal2 s 144816 0 144872 400 6 la_data_out[15]
port 214 nsew signal output
rlabel metal2 s 147504 0 147560 400 6 la_data_out[16]
port 215 nsew signal output
rlabel metal2 s 150192 0 150248 400 6 la_data_out[17]
port 216 nsew signal output
rlabel metal2 s 152880 0 152936 400 6 la_data_out[18]
port 217 nsew signal output
rlabel metal2 s 155568 0 155624 400 6 la_data_out[19]
port 218 nsew signal output
rlabel metal2 s 107184 0 107240 400 6 la_data_out[1]
port 219 nsew signal output
rlabel metal2 s 158256 0 158312 400 6 la_data_out[20]
port 220 nsew signal output
rlabel metal2 s 160944 0 161000 400 6 la_data_out[21]
port 221 nsew signal output
rlabel metal2 s 163632 0 163688 400 6 la_data_out[22]
port 222 nsew signal output
rlabel metal2 s 166320 0 166376 400 6 la_data_out[23]
port 223 nsew signal output
rlabel metal2 s 169008 0 169064 400 6 la_data_out[24]
port 224 nsew signal output
rlabel metal2 s 171696 0 171752 400 6 la_data_out[25]
port 225 nsew signal output
rlabel metal2 s 174384 0 174440 400 6 la_data_out[26]
port 226 nsew signal output
rlabel metal2 s 177072 0 177128 400 6 la_data_out[27]
port 227 nsew signal output
rlabel metal2 s 179760 0 179816 400 6 la_data_out[28]
port 228 nsew signal output
rlabel metal2 s 182448 0 182504 400 6 la_data_out[29]
port 229 nsew signal output
rlabel metal2 s 109872 0 109928 400 6 la_data_out[2]
port 230 nsew signal output
rlabel metal2 s 185136 0 185192 400 6 la_data_out[30]
port 231 nsew signal output
rlabel metal2 s 187824 0 187880 400 6 la_data_out[31]
port 232 nsew signal output
rlabel metal2 s 190512 0 190568 400 6 la_data_out[32]
port 233 nsew signal output
rlabel metal2 s 193200 0 193256 400 6 la_data_out[33]
port 234 nsew signal output
rlabel metal2 s 195888 0 195944 400 6 la_data_out[34]
port 235 nsew signal output
rlabel metal2 s 198576 0 198632 400 6 la_data_out[35]
port 236 nsew signal output
rlabel metal2 s 201264 0 201320 400 6 la_data_out[36]
port 237 nsew signal output
rlabel metal2 s 203952 0 204008 400 6 la_data_out[37]
port 238 nsew signal output
rlabel metal2 s 206640 0 206696 400 6 la_data_out[38]
port 239 nsew signal output
rlabel metal2 s 209328 0 209384 400 6 la_data_out[39]
port 240 nsew signal output
rlabel metal2 s 112560 0 112616 400 6 la_data_out[3]
port 241 nsew signal output
rlabel metal2 s 212016 0 212072 400 6 la_data_out[40]
port 242 nsew signal output
rlabel metal2 s 214704 0 214760 400 6 la_data_out[41]
port 243 nsew signal output
rlabel metal2 s 217392 0 217448 400 6 la_data_out[42]
port 244 nsew signal output
rlabel metal2 s 220080 0 220136 400 6 la_data_out[43]
port 245 nsew signal output
rlabel metal2 s 222768 0 222824 400 6 la_data_out[44]
port 246 nsew signal output
rlabel metal2 s 225456 0 225512 400 6 la_data_out[45]
port 247 nsew signal output
rlabel metal2 s 228144 0 228200 400 6 la_data_out[46]
port 248 nsew signal output
rlabel metal2 s 230832 0 230888 400 6 la_data_out[47]
port 249 nsew signal output
rlabel metal2 s 233520 0 233576 400 6 la_data_out[48]
port 250 nsew signal output
rlabel metal2 s 236208 0 236264 400 6 la_data_out[49]
port 251 nsew signal output
rlabel metal2 s 115248 0 115304 400 6 la_data_out[4]
port 252 nsew signal output
rlabel metal2 s 238896 0 238952 400 6 la_data_out[50]
port 253 nsew signal output
rlabel metal2 s 241584 0 241640 400 6 la_data_out[51]
port 254 nsew signal output
rlabel metal2 s 244272 0 244328 400 6 la_data_out[52]
port 255 nsew signal output
rlabel metal2 s 246960 0 247016 400 6 la_data_out[53]
port 256 nsew signal output
rlabel metal2 s 249648 0 249704 400 6 la_data_out[54]
port 257 nsew signal output
rlabel metal2 s 252336 0 252392 400 6 la_data_out[55]
port 258 nsew signal output
rlabel metal2 s 255024 0 255080 400 6 la_data_out[56]
port 259 nsew signal output
rlabel metal2 s 257712 0 257768 400 6 la_data_out[57]
port 260 nsew signal output
rlabel metal2 s 260400 0 260456 400 6 la_data_out[58]
port 261 nsew signal output
rlabel metal2 s 263088 0 263144 400 6 la_data_out[59]
port 262 nsew signal output
rlabel metal2 s 117936 0 117992 400 6 la_data_out[5]
port 263 nsew signal output
rlabel metal2 s 265776 0 265832 400 6 la_data_out[60]
port 264 nsew signal output
rlabel metal2 s 268464 0 268520 400 6 la_data_out[61]
port 265 nsew signal output
rlabel metal2 s 271152 0 271208 400 6 la_data_out[62]
port 266 nsew signal output
rlabel metal2 s 273840 0 273896 400 6 la_data_out[63]
port 267 nsew signal output
rlabel metal2 s 120624 0 120680 400 6 la_data_out[6]
port 268 nsew signal output
rlabel metal2 s 123312 0 123368 400 6 la_data_out[7]
port 269 nsew signal output
rlabel metal2 s 126000 0 126056 400 6 la_data_out[8]
port 270 nsew signal output
rlabel metal2 s 128688 0 128744 400 6 la_data_out[9]
port 271 nsew signal output
rlabel metal2 s 105392 0 105448 400 6 la_oenb[0]
port 272 nsew signal input
rlabel metal2 s 132272 0 132328 400 6 la_oenb[10]
port 273 nsew signal input
rlabel metal2 s 134960 0 135016 400 6 la_oenb[11]
port 274 nsew signal input
rlabel metal2 s 137648 0 137704 400 6 la_oenb[12]
port 275 nsew signal input
rlabel metal2 s 140336 0 140392 400 6 la_oenb[13]
port 276 nsew signal input
rlabel metal2 s 143024 0 143080 400 6 la_oenb[14]
port 277 nsew signal input
rlabel metal2 s 145712 0 145768 400 6 la_oenb[15]
port 278 nsew signal input
rlabel metal2 s 148400 0 148456 400 6 la_oenb[16]
port 279 nsew signal input
rlabel metal2 s 151088 0 151144 400 6 la_oenb[17]
port 280 nsew signal input
rlabel metal2 s 153776 0 153832 400 6 la_oenb[18]
port 281 nsew signal input
rlabel metal2 s 156464 0 156520 400 6 la_oenb[19]
port 282 nsew signal input
rlabel metal2 s 108080 0 108136 400 6 la_oenb[1]
port 283 nsew signal input
rlabel metal2 s 159152 0 159208 400 6 la_oenb[20]
port 284 nsew signal input
rlabel metal2 s 161840 0 161896 400 6 la_oenb[21]
port 285 nsew signal input
rlabel metal2 s 164528 0 164584 400 6 la_oenb[22]
port 286 nsew signal input
rlabel metal2 s 167216 0 167272 400 6 la_oenb[23]
port 287 nsew signal input
rlabel metal2 s 169904 0 169960 400 6 la_oenb[24]
port 288 nsew signal input
rlabel metal2 s 172592 0 172648 400 6 la_oenb[25]
port 289 nsew signal input
rlabel metal2 s 175280 0 175336 400 6 la_oenb[26]
port 290 nsew signal input
rlabel metal2 s 177968 0 178024 400 6 la_oenb[27]
port 291 nsew signal input
rlabel metal2 s 180656 0 180712 400 6 la_oenb[28]
port 292 nsew signal input
rlabel metal2 s 183344 0 183400 400 6 la_oenb[29]
port 293 nsew signal input
rlabel metal2 s 110768 0 110824 400 6 la_oenb[2]
port 294 nsew signal input
rlabel metal2 s 186032 0 186088 400 6 la_oenb[30]
port 295 nsew signal input
rlabel metal2 s 188720 0 188776 400 6 la_oenb[31]
port 296 nsew signal input
rlabel metal2 s 191408 0 191464 400 6 la_oenb[32]
port 297 nsew signal input
rlabel metal2 s 194096 0 194152 400 6 la_oenb[33]
port 298 nsew signal input
rlabel metal2 s 196784 0 196840 400 6 la_oenb[34]
port 299 nsew signal input
rlabel metal2 s 199472 0 199528 400 6 la_oenb[35]
port 300 nsew signal input
rlabel metal2 s 202160 0 202216 400 6 la_oenb[36]
port 301 nsew signal input
rlabel metal2 s 204848 0 204904 400 6 la_oenb[37]
port 302 nsew signal input
rlabel metal2 s 207536 0 207592 400 6 la_oenb[38]
port 303 nsew signal input
rlabel metal2 s 210224 0 210280 400 6 la_oenb[39]
port 304 nsew signal input
rlabel metal2 s 113456 0 113512 400 6 la_oenb[3]
port 305 nsew signal input
rlabel metal2 s 212912 0 212968 400 6 la_oenb[40]
port 306 nsew signal input
rlabel metal2 s 215600 0 215656 400 6 la_oenb[41]
port 307 nsew signal input
rlabel metal2 s 218288 0 218344 400 6 la_oenb[42]
port 308 nsew signal input
rlabel metal2 s 220976 0 221032 400 6 la_oenb[43]
port 309 nsew signal input
rlabel metal2 s 223664 0 223720 400 6 la_oenb[44]
port 310 nsew signal input
rlabel metal2 s 226352 0 226408 400 6 la_oenb[45]
port 311 nsew signal input
rlabel metal2 s 229040 0 229096 400 6 la_oenb[46]
port 312 nsew signal input
rlabel metal2 s 231728 0 231784 400 6 la_oenb[47]
port 313 nsew signal input
rlabel metal2 s 234416 0 234472 400 6 la_oenb[48]
port 314 nsew signal input
rlabel metal2 s 237104 0 237160 400 6 la_oenb[49]
port 315 nsew signal input
rlabel metal2 s 116144 0 116200 400 6 la_oenb[4]
port 316 nsew signal input
rlabel metal2 s 239792 0 239848 400 6 la_oenb[50]
port 317 nsew signal input
rlabel metal2 s 242480 0 242536 400 6 la_oenb[51]
port 318 nsew signal input
rlabel metal2 s 245168 0 245224 400 6 la_oenb[52]
port 319 nsew signal input
rlabel metal2 s 247856 0 247912 400 6 la_oenb[53]
port 320 nsew signal input
rlabel metal2 s 250544 0 250600 400 6 la_oenb[54]
port 321 nsew signal input
rlabel metal2 s 253232 0 253288 400 6 la_oenb[55]
port 322 nsew signal input
rlabel metal2 s 255920 0 255976 400 6 la_oenb[56]
port 323 nsew signal input
rlabel metal2 s 258608 0 258664 400 6 la_oenb[57]
port 324 nsew signal input
rlabel metal2 s 261296 0 261352 400 6 la_oenb[58]
port 325 nsew signal input
rlabel metal2 s 263984 0 264040 400 6 la_oenb[59]
port 326 nsew signal input
rlabel metal2 s 118832 0 118888 400 6 la_oenb[5]
port 327 nsew signal input
rlabel metal2 s 266672 0 266728 400 6 la_oenb[60]
port 328 nsew signal input
rlabel metal2 s 269360 0 269416 400 6 la_oenb[61]
port 329 nsew signal input
rlabel metal2 s 272048 0 272104 400 6 la_oenb[62]
port 330 nsew signal input
rlabel metal2 s 274736 0 274792 400 6 la_oenb[63]
port 331 nsew signal input
rlabel metal2 s 121520 0 121576 400 6 la_oenb[6]
port 332 nsew signal input
rlabel metal2 s 124208 0 124264 400 6 la_oenb[7]
port 333 nsew signal input
rlabel metal2 s 126896 0 126952 400 6 la_oenb[8]
port 334 nsew signal input
rlabel metal2 s 129584 0 129640 400 6 la_oenb[9]
port 335 nsew signal input
rlabel metal2 s 275632 0 275688 400 6 user_clock2
port 336 nsew signal input
rlabel metal2 s 276528 0 276584 400 6 user_irq[0]
port 337 nsew signal output
rlabel metal2 s 277424 0 277480 400 6 user_irq[1]
port 338 nsew signal output
rlabel metal2 s 278320 0 278376 400 6 user_irq[2]
port 339 nsew signal output
rlabel metal4 s 2224 1538 2384 286974 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 286974 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 286974 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 286974 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 286974 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 286974 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 286974 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 286974 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 286974 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 286974 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 286974 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 286974 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 286974 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 201904 1538 202064 286974 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 217264 1538 217424 286974 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 232624 1538 232784 286974 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 247984 1538 248144 286974 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 263344 1538 263504 286974 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 278704 1538 278864 286974 6 vdd
port 340 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 286974 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 286974 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 286974 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 286974 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 286974 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 286974 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 286974 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 286974 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 286974 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 286974 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 286974 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 286974 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 286974 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 209584 1538 209744 286974 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 224944 1538 225104 286974 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 240304 1538 240464 286974 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 255664 1538 255824 286974 6 vss
port 341 nsew ground bidirectional
rlabel metal4 s 271024 1538 271184 286974 6 vss
port 341 nsew ground bidirectional
rlabel metal2 s 8624 0 8680 400 6 wb_clk_i
port 342 nsew signal input
rlabel metal2 s 9520 0 9576 400 6 wb_rst_i
port 343 nsew signal input
rlabel metal2 s 10416 0 10472 400 6 wbs_ack_o
port 344 nsew signal output
rlabel metal2 s 14000 0 14056 400 6 wbs_adr_i[0]
port 345 nsew signal input
rlabel metal2 s 44464 0 44520 400 6 wbs_adr_i[10]
port 346 nsew signal input
rlabel metal2 s 47152 0 47208 400 6 wbs_adr_i[11]
port 347 nsew signal input
rlabel metal2 s 49840 0 49896 400 6 wbs_adr_i[12]
port 348 nsew signal input
rlabel metal2 s 52528 0 52584 400 6 wbs_adr_i[13]
port 349 nsew signal input
rlabel metal2 s 55216 0 55272 400 6 wbs_adr_i[14]
port 350 nsew signal input
rlabel metal2 s 57904 0 57960 400 6 wbs_adr_i[15]
port 351 nsew signal input
rlabel metal2 s 60592 0 60648 400 6 wbs_adr_i[16]
port 352 nsew signal input
rlabel metal2 s 63280 0 63336 400 6 wbs_adr_i[17]
port 353 nsew signal input
rlabel metal2 s 65968 0 66024 400 6 wbs_adr_i[18]
port 354 nsew signal input
rlabel metal2 s 68656 0 68712 400 6 wbs_adr_i[19]
port 355 nsew signal input
rlabel metal2 s 17584 0 17640 400 6 wbs_adr_i[1]
port 356 nsew signal input
rlabel metal2 s 71344 0 71400 400 6 wbs_adr_i[20]
port 357 nsew signal input
rlabel metal2 s 74032 0 74088 400 6 wbs_adr_i[21]
port 358 nsew signal input
rlabel metal2 s 76720 0 76776 400 6 wbs_adr_i[22]
port 359 nsew signal input
rlabel metal2 s 79408 0 79464 400 6 wbs_adr_i[23]
port 360 nsew signal input
rlabel metal2 s 82096 0 82152 400 6 wbs_adr_i[24]
port 361 nsew signal input
rlabel metal2 s 84784 0 84840 400 6 wbs_adr_i[25]
port 362 nsew signal input
rlabel metal2 s 87472 0 87528 400 6 wbs_adr_i[26]
port 363 nsew signal input
rlabel metal2 s 90160 0 90216 400 6 wbs_adr_i[27]
port 364 nsew signal input
rlabel metal2 s 92848 0 92904 400 6 wbs_adr_i[28]
port 365 nsew signal input
rlabel metal2 s 95536 0 95592 400 6 wbs_adr_i[29]
port 366 nsew signal input
rlabel metal2 s 21168 0 21224 400 6 wbs_adr_i[2]
port 367 nsew signal input
rlabel metal2 s 98224 0 98280 400 6 wbs_adr_i[30]
port 368 nsew signal input
rlabel metal2 s 100912 0 100968 400 6 wbs_adr_i[31]
port 369 nsew signal input
rlabel metal2 s 24752 0 24808 400 6 wbs_adr_i[3]
port 370 nsew signal input
rlabel metal2 s 28336 0 28392 400 6 wbs_adr_i[4]
port 371 nsew signal input
rlabel metal2 s 31024 0 31080 400 6 wbs_adr_i[5]
port 372 nsew signal input
rlabel metal2 s 33712 0 33768 400 6 wbs_adr_i[6]
port 373 nsew signal input
rlabel metal2 s 36400 0 36456 400 6 wbs_adr_i[7]
port 374 nsew signal input
rlabel metal2 s 39088 0 39144 400 6 wbs_adr_i[8]
port 375 nsew signal input
rlabel metal2 s 41776 0 41832 400 6 wbs_adr_i[9]
port 376 nsew signal input
rlabel metal2 s 11312 0 11368 400 6 wbs_cyc_i
port 377 nsew signal input
rlabel metal2 s 14896 0 14952 400 6 wbs_dat_i[0]
port 378 nsew signal input
rlabel metal2 s 45360 0 45416 400 6 wbs_dat_i[10]
port 379 nsew signal input
rlabel metal2 s 48048 0 48104 400 6 wbs_dat_i[11]
port 380 nsew signal input
rlabel metal2 s 50736 0 50792 400 6 wbs_dat_i[12]
port 381 nsew signal input
rlabel metal2 s 53424 0 53480 400 6 wbs_dat_i[13]
port 382 nsew signal input
rlabel metal2 s 56112 0 56168 400 6 wbs_dat_i[14]
port 383 nsew signal input
rlabel metal2 s 58800 0 58856 400 6 wbs_dat_i[15]
port 384 nsew signal input
rlabel metal2 s 61488 0 61544 400 6 wbs_dat_i[16]
port 385 nsew signal input
rlabel metal2 s 64176 0 64232 400 6 wbs_dat_i[17]
port 386 nsew signal input
rlabel metal2 s 66864 0 66920 400 6 wbs_dat_i[18]
port 387 nsew signal input
rlabel metal2 s 69552 0 69608 400 6 wbs_dat_i[19]
port 388 nsew signal input
rlabel metal2 s 18480 0 18536 400 6 wbs_dat_i[1]
port 389 nsew signal input
rlabel metal2 s 72240 0 72296 400 6 wbs_dat_i[20]
port 390 nsew signal input
rlabel metal2 s 74928 0 74984 400 6 wbs_dat_i[21]
port 391 nsew signal input
rlabel metal2 s 77616 0 77672 400 6 wbs_dat_i[22]
port 392 nsew signal input
rlabel metal2 s 80304 0 80360 400 6 wbs_dat_i[23]
port 393 nsew signal input
rlabel metal2 s 82992 0 83048 400 6 wbs_dat_i[24]
port 394 nsew signal input
rlabel metal2 s 85680 0 85736 400 6 wbs_dat_i[25]
port 395 nsew signal input
rlabel metal2 s 88368 0 88424 400 6 wbs_dat_i[26]
port 396 nsew signal input
rlabel metal2 s 91056 0 91112 400 6 wbs_dat_i[27]
port 397 nsew signal input
rlabel metal2 s 93744 0 93800 400 6 wbs_dat_i[28]
port 398 nsew signal input
rlabel metal2 s 96432 0 96488 400 6 wbs_dat_i[29]
port 399 nsew signal input
rlabel metal2 s 22064 0 22120 400 6 wbs_dat_i[2]
port 400 nsew signal input
rlabel metal2 s 99120 0 99176 400 6 wbs_dat_i[30]
port 401 nsew signal input
rlabel metal2 s 101808 0 101864 400 6 wbs_dat_i[31]
port 402 nsew signal input
rlabel metal2 s 25648 0 25704 400 6 wbs_dat_i[3]
port 403 nsew signal input
rlabel metal2 s 29232 0 29288 400 6 wbs_dat_i[4]
port 404 nsew signal input
rlabel metal2 s 31920 0 31976 400 6 wbs_dat_i[5]
port 405 nsew signal input
rlabel metal2 s 34608 0 34664 400 6 wbs_dat_i[6]
port 406 nsew signal input
rlabel metal2 s 37296 0 37352 400 6 wbs_dat_i[7]
port 407 nsew signal input
rlabel metal2 s 39984 0 40040 400 6 wbs_dat_i[8]
port 408 nsew signal input
rlabel metal2 s 42672 0 42728 400 6 wbs_dat_i[9]
port 409 nsew signal input
rlabel metal2 s 15792 0 15848 400 6 wbs_dat_o[0]
port 410 nsew signal output
rlabel metal2 s 46256 0 46312 400 6 wbs_dat_o[10]
port 411 nsew signal output
rlabel metal2 s 48944 0 49000 400 6 wbs_dat_o[11]
port 412 nsew signal output
rlabel metal2 s 51632 0 51688 400 6 wbs_dat_o[12]
port 413 nsew signal output
rlabel metal2 s 54320 0 54376 400 6 wbs_dat_o[13]
port 414 nsew signal output
rlabel metal2 s 57008 0 57064 400 6 wbs_dat_o[14]
port 415 nsew signal output
rlabel metal2 s 59696 0 59752 400 6 wbs_dat_o[15]
port 416 nsew signal output
rlabel metal2 s 62384 0 62440 400 6 wbs_dat_o[16]
port 417 nsew signal output
rlabel metal2 s 65072 0 65128 400 6 wbs_dat_o[17]
port 418 nsew signal output
rlabel metal2 s 67760 0 67816 400 6 wbs_dat_o[18]
port 419 nsew signal output
rlabel metal2 s 70448 0 70504 400 6 wbs_dat_o[19]
port 420 nsew signal output
rlabel metal2 s 19376 0 19432 400 6 wbs_dat_o[1]
port 421 nsew signal output
rlabel metal2 s 73136 0 73192 400 6 wbs_dat_o[20]
port 422 nsew signal output
rlabel metal2 s 75824 0 75880 400 6 wbs_dat_o[21]
port 423 nsew signal output
rlabel metal2 s 78512 0 78568 400 6 wbs_dat_o[22]
port 424 nsew signal output
rlabel metal2 s 81200 0 81256 400 6 wbs_dat_o[23]
port 425 nsew signal output
rlabel metal2 s 83888 0 83944 400 6 wbs_dat_o[24]
port 426 nsew signal output
rlabel metal2 s 86576 0 86632 400 6 wbs_dat_o[25]
port 427 nsew signal output
rlabel metal2 s 89264 0 89320 400 6 wbs_dat_o[26]
port 428 nsew signal output
rlabel metal2 s 91952 0 92008 400 6 wbs_dat_o[27]
port 429 nsew signal output
rlabel metal2 s 94640 0 94696 400 6 wbs_dat_o[28]
port 430 nsew signal output
rlabel metal2 s 97328 0 97384 400 6 wbs_dat_o[29]
port 431 nsew signal output
rlabel metal2 s 22960 0 23016 400 6 wbs_dat_o[2]
port 432 nsew signal output
rlabel metal2 s 100016 0 100072 400 6 wbs_dat_o[30]
port 433 nsew signal output
rlabel metal2 s 102704 0 102760 400 6 wbs_dat_o[31]
port 434 nsew signal output
rlabel metal2 s 26544 0 26600 400 6 wbs_dat_o[3]
port 435 nsew signal output
rlabel metal2 s 30128 0 30184 400 6 wbs_dat_o[4]
port 436 nsew signal output
rlabel metal2 s 32816 0 32872 400 6 wbs_dat_o[5]
port 437 nsew signal output
rlabel metal2 s 35504 0 35560 400 6 wbs_dat_o[6]
port 438 nsew signal output
rlabel metal2 s 38192 0 38248 400 6 wbs_dat_o[7]
port 439 nsew signal output
rlabel metal2 s 40880 0 40936 400 6 wbs_dat_o[8]
port 440 nsew signal output
rlabel metal2 s 43568 0 43624 400 6 wbs_dat_o[9]
port 441 nsew signal output
rlabel metal2 s 16688 0 16744 400 6 wbs_sel_i[0]
port 442 nsew signal input
rlabel metal2 s 20272 0 20328 400 6 wbs_sel_i[1]
port 443 nsew signal input
rlabel metal2 s 23856 0 23912 400 6 wbs_sel_i[2]
port 444 nsew signal input
rlabel metal2 s 27440 0 27496 400 6 wbs_sel_i[3]
port 445 nsew signal input
rlabel metal2 s 12208 0 12264 400 6 wbs_stb_i
port 446 nsew signal input
rlabel metal2 s 13104 0 13160 400 6 wbs_we_i
port 447 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 287047 288839
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 243591442
string GDS_FILE /mnt/r/work/Rift2Go_2300_GF180_MPW1_1/openlane/user_proj_example/runs/23_11_02_09_53/results/signoff/rift2Wrap.magic.gds
string GDS_START 731710
<< end >>

