VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO rift2Wrap
  CLASS BLOCK ;
  FOREIGN rift2Wrap ;
  ORIGIN 0.000 0.000 ;
  SIZE 2870.470 BY 2888.390 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 1174.880 2870.470 1175.440 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2189.600 2884.390 2190.160 2888.390 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1871.520 2884.390 1872.080 2888.390 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1553.440 2884.390 1554.000 2888.390 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1235.360 2884.390 1235.920 2888.390 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 917.280 2884.390 917.840 2888.390 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 599.200 2884.390 599.760 2888.390 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 281.120 2884.390 281.680 2888.390 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2838.080 4.000 2838.640 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2627.520 4.000 2628.080 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2416.960 4.000 2417.520 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 1389.920 2870.470 1390.480 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2206.400 4.000 2206.960 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1995.840 4.000 1996.400 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1785.280 4.000 1785.840 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1574.720 4.000 1575.280 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1364.160 4.000 1364.720 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1153.600 4.000 1154.160 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 943.040 4.000 943.600 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 732.480 4.000 733.040 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 521.920 4.000 522.480 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 1604.960 2870.470 1605.520 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 1820.000 2870.470 1820.560 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 2035.040 2870.470 2035.600 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 2250.080 2870.470 2250.640 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 2465.120 2870.470 2465.680 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 2680.160 2870.470 2680.720 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2825.760 2884.390 2826.320 2888.390 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2507.680 2884.390 2508.240 2888.390 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 45.920 2870.470 46.480 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 1873.760 2870.470 1874.320 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 2088.800 2870.470 2089.360 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 2303.840 2870.470 2304.400 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 2518.880 2870.470 2519.440 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 2733.920 2870.470 2734.480 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2746.240 2884.390 2746.800 2888.390 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2428.160 2884.390 2428.720 2888.390 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2110.080 2884.390 2110.640 2888.390 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1792.000 2884.390 1792.560 2888.390 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1473.920 2884.390 1474.480 2888.390 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 207.200 2870.470 207.760 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1155.840 2884.390 1156.400 2888.390 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 837.760 2884.390 838.320 2888.390 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.369000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 519.680 2884.390 520.240 2888.390 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.408000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 201.600 2884.390 202.160 2888.390 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.612000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2785.440 4.000 2786.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2574.880 4.000 2575.440 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2364.320 4.000 2364.880 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2153.760 4.000 2154.320 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1943.200 4.000 1943.760 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1732.640 4.000 1733.200 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 368.480 2870.470 369.040 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1522.080 4.000 1522.640 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1311.520 4.000 1312.080 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1100.960 4.000 1101.520 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 890.400 4.000 890.960 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 679.840 4.000 680.400 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 469.280 4.000 469.840 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 311.360 4.000 311.920 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 153.440 4.000 154.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 529.760 2870.470 530.320 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 691.040 2870.470 691.600 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 852.320 2870.470 852.880 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 1013.600 2870.470 1014.160 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 1228.640 2870.470 1229.200 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 1443.680 2870.470 1444.240 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 1658.720 2870.470 1659.280 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 153.440 2870.470 154.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 1981.280 2870.470 1981.840 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 2196.320 2870.470 2196.880 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 2411.360 2870.470 2411.920 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 2626.400 2870.470 2626.960 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 2841.440 2870.470 2842.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2587.200 2884.390 2587.760 2888.390 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2269.120 2884.390 2269.680 2888.390 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1951.040 2884.390 1951.600 2888.390 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1632.960 2884.390 1633.520 2888.390 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1314.880 2884.390 1315.440 2888.390 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 314.720 2870.470 315.280 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 996.800 2884.390 997.360 2888.390 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 2884.390 679.280 2888.390 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 360.640 2884.390 361.200 2888.390 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 42.560 2884.390 43.120 2888.390 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2680.160 4.000 2680.720 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2469.600 4.000 2470.160 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2259.040 4.000 2259.600 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2048.480 4.000 2049.040 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1837.920 4.000 1838.480 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1627.360 4.000 1627.920 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 476.000 2870.470 476.560 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1416.800 4.000 1417.360 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1206.240 4.000 1206.800 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 995.680 4.000 996.240 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 785.120 4.000 785.680 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 574.560 4.000 575.120 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 364.000 4.000 364.560 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 206.080 4.000 206.640 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 48.160 4.000 48.720 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 637.280 2870.470 637.840 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 798.560 2870.470 799.120 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 959.840 2870.470 960.400 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 1121.120 2870.470 1121.680 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 1336.160 2870.470 1336.720 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 1551.200 2870.470 1551.760 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 1766.240 2870.470 1766.800 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 99.680 2870.470 100.240 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 1927.520 2870.470 1928.080 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 2142.560 2870.470 2143.120 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 2357.600 2870.470 2358.160 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 2572.640 2870.470 2573.200 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 2787.680 2870.470 2788.240 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2666.720 2884.390 2667.280 2888.390 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2348.640 2884.390 2349.200 2888.390 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 2030.560 2884.390 2031.120 2888.390 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1712.480 2884.390 1713.040 2888.390 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1394.400 2884.390 1394.960 2888.390 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 260.960 2870.470 261.520 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1076.320 2884.390 1076.880 2888.390 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 758.240 2884.390 758.800 2888.390 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 440.160 2884.390 440.720 2888.390 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 122.080 2884.390 122.640 2888.390 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2732.800 4.000 2733.360 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2522.240 4.000 2522.800 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2311.680 4.000 2312.240 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 2101.120 4.000 2101.680 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1890.560 4.000 1891.120 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1680.000 4.000 1680.560 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 422.240 2870.470 422.800 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1469.440 4.000 1470.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1258.880 4.000 1259.440 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 1048.320 4.000 1048.880 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 837.760 4.000 838.320 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 627.200 4.000 627.760 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 416.640 4.000 417.200 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 258.720 4.000 259.280 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 100.800 4.000 101.360 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 583.520 2870.470 584.080 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 744.800 2870.470 745.360 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 906.080 2870.470 906.640 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 1067.360 2870.470 1067.920 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 1282.400 2870.470 1282.960 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 1497.440 2870.470 1498.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 2866.470 1712.480 2870.470 1713.040 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1036.000 0.000 1036.560 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1304.800 0.000 1305.360 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1331.680 0.000 1332.240 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1358.560 0.000 1359.120 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1385.440 0.000 1386.000 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1412.320 0.000 1412.880 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1439.200 0.000 1439.760 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1466.080 0.000 1466.640 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1492.960 0.000 1493.520 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1519.840 0.000 1520.400 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1546.720 0.000 1547.280 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1062.880 0.000 1063.440 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1573.600 0.000 1574.160 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1600.480 0.000 1601.040 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1627.360 0.000 1627.920 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1654.240 0.000 1654.800 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1681.120 0.000 1681.680 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1708.000 0.000 1708.560 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1734.880 0.000 1735.440 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1761.760 0.000 1762.320 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1788.640 0.000 1789.200 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1815.520 0.000 1816.080 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1089.760 0.000 1090.320 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1842.400 0.000 1842.960 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1869.280 0.000 1869.840 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1896.160 0.000 1896.720 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1923.040 0.000 1923.600 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1949.920 0.000 1950.480 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1976.800 0.000 1977.360 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2003.680 0.000 2004.240 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2030.560 0.000 2031.120 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2057.440 0.000 2058.000 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2084.320 0.000 2084.880 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1116.640 0.000 1117.200 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2111.200 0.000 2111.760 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2138.080 0.000 2138.640 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2164.960 0.000 2165.520 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2191.840 0.000 2192.400 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2218.720 0.000 2219.280 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2245.600 0.000 2246.160 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2272.480 0.000 2273.040 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2299.360 0.000 2299.920 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2326.240 0.000 2326.800 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2353.120 0.000 2353.680 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1143.520 0.000 1144.080 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2380.000 0.000 2380.560 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2406.880 0.000 2407.440 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2433.760 0.000 2434.320 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2460.640 0.000 2461.200 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2487.520 0.000 2488.080 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2514.400 0.000 2514.960 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2541.280 0.000 2541.840 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2568.160 0.000 2568.720 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2595.040 0.000 2595.600 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2621.920 0.000 2622.480 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1170.400 0.000 1170.960 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2648.800 0.000 2649.360 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2675.680 0.000 2676.240 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2702.560 0.000 2703.120 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2729.440 0.000 2730.000 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1197.280 0.000 1197.840 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1224.160 0.000 1224.720 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1251.040 0.000 1251.600 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1277.920 0.000 1278.480 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1044.960 0.000 1045.520 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1313.760 0.000 1314.320 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1340.640 0.000 1341.200 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1367.520 0.000 1368.080 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1394.400 0.000 1394.960 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1421.280 0.000 1421.840 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1448.160 0.000 1448.720 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1475.040 0.000 1475.600 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1501.920 0.000 1502.480 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1528.800 0.000 1529.360 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1555.680 0.000 1556.240 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1071.840 0.000 1072.400 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1582.560 0.000 1583.120 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1609.440 0.000 1610.000 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1636.320 0.000 1636.880 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1663.200 0.000 1663.760 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1690.080 0.000 1690.640 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1716.960 0.000 1717.520 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1743.840 0.000 1744.400 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1770.720 0.000 1771.280 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1797.600 0.000 1798.160 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1824.480 0.000 1825.040 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1098.720 0.000 1099.280 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1851.360 0.000 1851.920 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1878.240 0.000 1878.800 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1905.120 0.000 1905.680 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1932.000 0.000 1932.560 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1958.880 0.000 1959.440 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1985.760 0.000 1986.320 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2012.640 0.000 2013.200 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2039.520 0.000 2040.080 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2066.400 0.000 2066.960 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2093.280 0.000 2093.840 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1125.600 0.000 1126.160 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2120.160 0.000 2120.720 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2147.040 0.000 2147.600 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2173.920 0.000 2174.480 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2200.800 0.000 2201.360 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2227.680 0.000 2228.240 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2254.560 0.000 2255.120 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2281.440 0.000 2282.000 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2308.320 0.000 2308.880 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2335.200 0.000 2335.760 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2362.080 0.000 2362.640 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1152.480 0.000 1153.040 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2388.960 0.000 2389.520 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2415.840 0.000 2416.400 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2442.720 0.000 2443.280 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2469.600 0.000 2470.160 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2496.480 0.000 2497.040 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2523.360 0.000 2523.920 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2550.240 0.000 2550.800 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2577.120 0.000 2577.680 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2604.000 0.000 2604.560 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2630.880 0.000 2631.440 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1179.360 0.000 1179.920 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2657.760 0.000 2658.320 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2684.640 0.000 2685.200 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2711.520 0.000 2712.080 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2738.400 0.000 2738.960 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1206.240 0.000 1206.800 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1233.120 0.000 1233.680 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1260.000 0.000 1260.560 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1286.880 0.000 1287.440 4.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1053.920 0.000 1054.480 4.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1322.720 0.000 1323.280 4.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1349.600 0.000 1350.160 4.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1376.480 0.000 1377.040 4.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1403.360 0.000 1403.920 4.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1430.240 0.000 1430.800 4.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1457.120 0.000 1457.680 4.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1484.000 0.000 1484.560 4.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1510.880 0.000 1511.440 4.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1537.760 0.000 1538.320 4.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1564.640 0.000 1565.200 4.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1080.800 0.000 1081.360 4.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1591.520 0.000 1592.080 4.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1618.400 0.000 1618.960 4.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1645.280 0.000 1645.840 4.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1672.160 0.000 1672.720 4.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1699.040 0.000 1699.600 4.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1725.920 0.000 1726.480 4.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1752.800 0.000 1753.360 4.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1779.680 0.000 1780.240 4.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1806.560 0.000 1807.120 4.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1833.440 0.000 1834.000 4.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1107.680 0.000 1108.240 4.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1860.320 0.000 1860.880 4.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1887.200 0.000 1887.760 4.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1914.080 0.000 1914.640 4.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1940.960 0.000 1941.520 4.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1967.840 0.000 1968.400 4.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1994.720 0.000 1995.280 4.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2021.600 0.000 2022.160 4.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2048.480 0.000 2049.040 4.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2075.360 0.000 2075.920 4.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2102.240 0.000 2102.800 4.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1134.560 0.000 1135.120 4.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2129.120 0.000 2129.680 4.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2156.000 0.000 2156.560 4.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2182.880 0.000 2183.440 4.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2209.760 0.000 2210.320 4.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2236.640 0.000 2237.200 4.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2263.520 0.000 2264.080 4.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2290.400 0.000 2290.960 4.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2317.280 0.000 2317.840 4.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2344.160 0.000 2344.720 4.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2371.040 0.000 2371.600 4.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1161.440 0.000 1162.000 4.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2397.920 0.000 2398.480 4.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2424.800 0.000 2425.360 4.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2451.680 0.000 2452.240 4.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2478.560 0.000 2479.120 4.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2505.440 0.000 2506.000 4.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2532.320 0.000 2532.880 4.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2559.200 0.000 2559.760 4.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2586.080 0.000 2586.640 4.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2612.960 0.000 2613.520 4.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2639.840 0.000 2640.400 4.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1188.320 0.000 1188.880 4.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2666.720 0.000 2667.280 4.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2693.600 0.000 2694.160 4.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2720.480 0.000 2721.040 4.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 2747.360 0.000 2747.920 4.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1215.200 0.000 1215.760 4.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1242.080 0.000 1242.640 4.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1268.960 0.000 1269.520 4.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1295.840 0.000 1296.400 4.000 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 2756.320 0.000 2756.880 4.000 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2765.280 0.000 2765.840 4.000 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2774.240 0.000 2774.800 4.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 2783.200 0.000 2783.760 4.000 ;
    END
  END user_irq[2]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1097.440 15.380 1099.040 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1251.040 15.380 1252.640 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1404.640 15.380 1406.240 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1558.240 15.380 1559.840 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1711.840 15.380 1713.440 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1865.440 15.380 1867.040 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2019.040 15.380 2020.640 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2172.640 15.380 2174.240 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2326.240 15.380 2327.840 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2479.840 15.380 2481.440 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2633.440 15.380 2635.040 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2787.040 15.380 2788.640 2869.740 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1174.240 15.380 1175.840 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1327.840 15.380 1329.440 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1481.440 15.380 1483.040 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1635.040 15.380 1636.640 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1788.640 15.380 1790.240 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1942.240 15.380 1943.840 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2095.840 15.380 2097.440 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2249.440 15.380 2251.040 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2403.040 15.380 2404.640 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2556.640 15.380 2558.240 2869.740 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 2710.240 15.380 2711.840 2869.740 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 86.240 0.000 86.800 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 95.200 0.000 95.760 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 0.000 104.720 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 140.000 0.000 140.560 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 444.640 0.000 445.200 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 471.520 0.000 472.080 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 498.400 0.000 498.960 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 525.280 0.000 525.840 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 552.160 0.000 552.720 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 579.040 0.000 579.600 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 605.920 0.000 606.480 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 632.800 0.000 633.360 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 659.680 0.000 660.240 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 686.560 0.000 687.120 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 175.840 0.000 176.400 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 713.440 0.000 714.000 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 740.320 0.000 740.880 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 767.200 0.000 767.760 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 794.080 0.000 794.640 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 820.960 0.000 821.520 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 847.840 0.000 848.400 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 874.720 0.000 875.280 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 901.600 0.000 902.160 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 928.480 0.000 929.040 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 955.360 0.000 955.920 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 211.680 0.000 212.240 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 982.240 0.000 982.800 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1009.120 0.000 1009.680 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 247.520 0.000 248.080 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 283.360 0.000 283.920 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 310.240 0.000 310.800 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 337.120 0.000 337.680 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 364.000 0.000 364.560 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 390.880 0.000 391.440 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 417.760 0.000 418.320 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 113.120 0.000 113.680 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 148.960 0.000 149.520 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 453.600 0.000 454.160 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 480.480 0.000 481.040 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 507.360 0.000 507.920 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 534.240 0.000 534.800 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 561.120 0.000 561.680 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 588.000 0.000 588.560 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 614.880 0.000 615.440 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 641.760 0.000 642.320 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 668.640 0.000 669.200 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 695.520 0.000 696.080 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 184.800 0.000 185.360 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 722.400 0.000 722.960 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 749.280 0.000 749.840 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 776.160 0.000 776.720 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 803.040 0.000 803.600 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 829.920 0.000 830.480 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 856.800 0.000 857.360 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 883.680 0.000 884.240 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 910.560 0.000 911.120 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 937.440 0.000 938.000 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 964.320 0.000 964.880 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 220.640 0.000 221.200 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 991.200 0.000 991.760 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1018.080 0.000 1018.640 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 256.480 0.000 257.040 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 292.320 0.000 292.880 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 319.200 0.000 319.760 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 346.080 0.000 346.640 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 372.960 0.000 373.520 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 399.840 0.000 400.400 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 426.720 0.000 427.280 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 157.920 0.000 158.480 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 462.560 0.000 463.120 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 489.440 0.000 490.000 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 516.320 0.000 516.880 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 543.200 0.000 543.760 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 570.080 0.000 570.640 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 596.960 0.000 597.520 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 623.840 0.000 624.400 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 650.720 0.000 651.280 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 677.600 0.000 678.160 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 704.480 0.000 705.040 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 193.760 0.000 194.320 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 731.360 0.000 731.920 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 758.240 0.000 758.800 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 785.120 0.000 785.680 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 812.000 0.000 812.560 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 838.880 0.000 839.440 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 865.760 0.000 866.320 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 892.640 0.000 893.200 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 919.520 0.000 920.080 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 946.400 0.000 946.960 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 973.280 0.000 973.840 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 229.600 0.000 230.160 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1000.160 0.000 1000.720 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 1027.040 0.000 1027.600 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 265.440 0.000 266.000 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 301.280 0.000 301.840 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 328.160 0.000 328.720 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 355.040 0.000 355.600 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 381.920 0.000 382.480 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 408.800 0.000 409.360 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 435.680 0.000 436.240 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 166.880 0.000 167.440 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 202.720 0.000 203.280 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 238.560 0.000 239.120 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 274.400 0.000 274.960 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 122.080 0.000 122.640 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 131.040 0.000 131.600 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 8.550 2863.280 2872.650 ;
      LAYER Metal2 ;
        RECT 4.620 2884.090 42.260 2884.390 ;
        RECT 43.420 2884.090 121.780 2884.390 ;
        RECT 122.940 2884.090 201.300 2884.390 ;
        RECT 202.460 2884.090 280.820 2884.390 ;
        RECT 281.980 2884.090 360.340 2884.390 ;
        RECT 361.500 2884.090 439.860 2884.390 ;
        RECT 441.020 2884.090 519.380 2884.390 ;
        RECT 520.540 2884.090 598.900 2884.390 ;
        RECT 600.060 2884.090 678.420 2884.390 ;
        RECT 679.580 2884.090 757.940 2884.390 ;
        RECT 759.100 2884.090 837.460 2884.390 ;
        RECT 838.620 2884.090 916.980 2884.390 ;
        RECT 918.140 2884.090 996.500 2884.390 ;
        RECT 997.660 2884.090 1076.020 2884.390 ;
        RECT 1077.180 2884.090 1155.540 2884.390 ;
        RECT 1156.700 2884.090 1235.060 2884.390 ;
        RECT 1236.220 2884.090 1314.580 2884.390 ;
        RECT 1315.740 2884.090 1394.100 2884.390 ;
        RECT 1395.260 2884.090 1473.620 2884.390 ;
        RECT 1474.780 2884.090 1553.140 2884.390 ;
        RECT 1554.300 2884.090 1632.660 2884.390 ;
        RECT 1633.820 2884.090 1712.180 2884.390 ;
        RECT 1713.340 2884.090 1791.700 2884.390 ;
        RECT 1792.860 2884.090 1871.220 2884.390 ;
        RECT 1872.380 2884.090 1950.740 2884.390 ;
        RECT 1951.900 2884.090 2030.260 2884.390 ;
        RECT 2031.420 2884.090 2109.780 2884.390 ;
        RECT 2110.940 2884.090 2189.300 2884.390 ;
        RECT 2190.460 2884.090 2268.820 2884.390 ;
        RECT 2269.980 2884.090 2348.340 2884.390 ;
        RECT 2349.500 2884.090 2427.860 2884.390 ;
        RECT 2429.020 2884.090 2507.380 2884.390 ;
        RECT 2508.540 2884.090 2586.900 2884.390 ;
        RECT 2588.060 2884.090 2666.420 2884.390 ;
        RECT 2667.580 2884.090 2745.940 2884.390 ;
        RECT 2747.100 2884.090 2825.460 2884.390 ;
        RECT 2826.620 2884.090 2863.700 2884.390 ;
        RECT 4.620 4.300 2863.700 2884.090 ;
        RECT 4.620 2.890 85.940 4.300 ;
        RECT 87.100 2.890 94.900 4.300 ;
        RECT 96.060 2.890 103.860 4.300 ;
        RECT 105.020 2.890 112.820 4.300 ;
        RECT 113.980 2.890 121.780 4.300 ;
        RECT 122.940 2.890 130.740 4.300 ;
        RECT 131.900 2.890 139.700 4.300 ;
        RECT 140.860 2.890 148.660 4.300 ;
        RECT 149.820 2.890 157.620 4.300 ;
        RECT 158.780 2.890 166.580 4.300 ;
        RECT 167.740 2.890 175.540 4.300 ;
        RECT 176.700 2.890 184.500 4.300 ;
        RECT 185.660 2.890 193.460 4.300 ;
        RECT 194.620 2.890 202.420 4.300 ;
        RECT 203.580 2.890 211.380 4.300 ;
        RECT 212.540 2.890 220.340 4.300 ;
        RECT 221.500 2.890 229.300 4.300 ;
        RECT 230.460 2.890 238.260 4.300 ;
        RECT 239.420 2.890 247.220 4.300 ;
        RECT 248.380 2.890 256.180 4.300 ;
        RECT 257.340 2.890 265.140 4.300 ;
        RECT 266.300 2.890 274.100 4.300 ;
        RECT 275.260 2.890 283.060 4.300 ;
        RECT 284.220 2.890 292.020 4.300 ;
        RECT 293.180 2.890 300.980 4.300 ;
        RECT 302.140 2.890 309.940 4.300 ;
        RECT 311.100 2.890 318.900 4.300 ;
        RECT 320.060 2.890 327.860 4.300 ;
        RECT 329.020 2.890 336.820 4.300 ;
        RECT 337.980 2.890 345.780 4.300 ;
        RECT 346.940 2.890 354.740 4.300 ;
        RECT 355.900 2.890 363.700 4.300 ;
        RECT 364.860 2.890 372.660 4.300 ;
        RECT 373.820 2.890 381.620 4.300 ;
        RECT 382.780 2.890 390.580 4.300 ;
        RECT 391.740 2.890 399.540 4.300 ;
        RECT 400.700 2.890 408.500 4.300 ;
        RECT 409.660 2.890 417.460 4.300 ;
        RECT 418.620 2.890 426.420 4.300 ;
        RECT 427.580 2.890 435.380 4.300 ;
        RECT 436.540 2.890 444.340 4.300 ;
        RECT 445.500 2.890 453.300 4.300 ;
        RECT 454.460 2.890 462.260 4.300 ;
        RECT 463.420 2.890 471.220 4.300 ;
        RECT 472.380 2.890 480.180 4.300 ;
        RECT 481.340 2.890 489.140 4.300 ;
        RECT 490.300 2.890 498.100 4.300 ;
        RECT 499.260 2.890 507.060 4.300 ;
        RECT 508.220 2.890 516.020 4.300 ;
        RECT 517.180 2.890 524.980 4.300 ;
        RECT 526.140 2.890 533.940 4.300 ;
        RECT 535.100 2.890 542.900 4.300 ;
        RECT 544.060 2.890 551.860 4.300 ;
        RECT 553.020 2.890 560.820 4.300 ;
        RECT 561.980 2.890 569.780 4.300 ;
        RECT 570.940 2.890 578.740 4.300 ;
        RECT 579.900 2.890 587.700 4.300 ;
        RECT 588.860 2.890 596.660 4.300 ;
        RECT 597.820 2.890 605.620 4.300 ;
        RECT 606.780 2.890 614.580 4.300 ;
        RECT 615.740 2.890 623.540 4.300 ;
        RECT 624.700 2.890 632.500 4.300 ;
        RECT 633.660 2.890 641.460 4.300 ;
        RECT 642.620 2.890 650.420 4.300 ;
        RECT 651.580 2.890 659.380 4.300 ;
        RECT 660.540 2.890 668.340 4.300 ;
        RECT 669.500 2.890 677.300 4.300 ;
        RECT 678.460 2.890 686.260 4.300 ;
        RECT 687.420 2.890 695.220 4.300 ;
        RECT 696.380 2.890 704.180 4.300 ;
        RECT 705.340 2.890 713.140 4.300 ;
        RECT 714.300 2.890 722.100 4.300 ;
        RECT 723.260 2.890 731.060 4.300 ;
        RECT 732.220 2.890 740.020 4.300 ;
        RECT 741.180 2.890 748.980 4.300 ;
        RECT 750.140 2.890 757.940 4.300 ;
        RECT 759.100 2.890 766.900 4.300 ;
        RECT 768.060 2.890 775.860 4.300 ;
        RECT 777.020 2.890 784.820 4.300 ;
        RECT 785.980 2.890 793.780 4.300 ;
        RECT 794.940 2.890 802.740 4.300 ;
        RECT 803.900 2.890 811.700 4.300 ;
        RECT 812.860 2.890 820.660 4.300 ;
        RECT 821.820 2.890 829.620 4.300 ;
        RECT 830.780 2.890 838.580 4.300 ;
        RECT 839.740 2.890 847.540 4.300 ;
        RECT 848.700 2.890 856.500 4.300 ;
        RECT 857.660 2.890 865.460 4.300 ;
        RECT 866.620 2.890 874.420 4.300 ;
        RECT 875.580 2.890 883.380 4.300 ;
        RECT 884.540 2.890 892.340 4.300 ;
        RECT 893.500 2.890 901.300 4.300 ;
        RECT 902.460 2.890 910.260 4.300 ;
        RECT 911.420 2.890 919.220 4.300 ;
        RECT 920.380 2.890 928.180 4.300 ;
        RECT 929.340 2.890 937.140 4.300 ;
        RECT 938.300 2.890 946.100 4.300 ;
        RECT 947.260 2.890 955.060 4.300 ;
        RECT 956.220 2.890 964.020 4.300 ;
        RECT 965.180 2.890 972.980 4.300 ;
        RECT 974.140 2.890 981.940 4.300 ;
        RECT 983.100 2.890 990.900 4.300 ;
        RECT 992.060 2.890 999.860 4.300 ;
        RECT 1001.020 2.890 1008.820 4.300 ;
        RECT 1009.980 2.890 1017.780 4.300 ;
        RECT 1018.940 2.890 1026.740 4.300 ;
        RECT 1027.900 2.890 1035.700 4.300 ;
        RECT 1036.860 2.890 1044.660 4.300 ;
        RECT 1045.820 2.890 1053.620 4.300 ;
        RECT 1054.780 2.890 1062.580 4.300 ;
        RECT 1063.740 2.890 1071.540 4.300 ;
        RECT 1072.700 2.890 1080.500 4.300 ;
        RECT 1081.660 2.890 1089.460 4.300 ;
        RECT 1090.620 2.890 1098.420 4.300 ;
        RECT 1099.580 2.890 1107.380 4.300 ;
        RECT 1108.540 2.890 1116.340 4.300 ;
        RECT 1117.500 2.890 1125.300 4.300 ;
        RECT 1126.460 2.890 1134.260 4.300 ;
        RECT 1135.420 2.890 1143.220 4.300 ;
        RECT 1144.380 2.890 1152.180 4.300 ;
        RECT 1153.340 2.890 1161.140 4.300 ;
        RECT 1162.300 2.890 1170.100 4.300 ;
        RECT 1171.260 2.890 1179.060 4.300 ;
        RECT 1180.220 2.890 1188.020 4.300 ;
        RECT 1189.180 2.890 1196.980 4.300 ;
        RECT 1198.140 2.890 1205.940 4.300 ;
        RECT 1207.100 2.890 1214.900 4.300 ;
        RECT 1216.060 2.890 1223.860 4.300 ;
        RECT 1225.020 2.890 1232.820 4.300 ;
        RECT 1233.980 2.890 1241.780 4.300 ;
        RECT 1242.940 2.890 1250.740 4.300 ;
        RECT 1251.900 2.890 1259.700 4.300 ;
        RECT 1260.860 2.890 1268.660 4.300 ;
        RECT 1269.820 2.890 1277.620 4.300 ;
        RECT 1278.780 2.890 1286.580 4.300 ;
        RECT 1287.740 2.890 1295.540 4.300 ;
        RECT 1296.700 2.890 1304.500 4.300 ;
        RECT 1305.660 2.890 1313.460 4.300 ;
        RECT 1314.620 2.890 1322.420 4.300 ;
        RECT 1323.580 2.890 1331.380 4.300 ;
        RECT 1332.540 2.890 1340.340 4.300 ;
        RECT 1341.500 2.890 1349.300 4.300 ;
        RECT 1350.460 2.890 1358.260 4.300 ;
        RECT 1359.420 2.890 1367.220 4.300 ;
        RECT 1368.380 2.890 1376.180 4.300 ;
        RECT 1377.340 2.890 1385.140 4.300 ;
        RECT 1386.300 2.890 1394.100 4.300 ;
        RECT 1395.260 2.890 1403.060 4.300 ;
        RECT 1404.220 2.890 1412.020 4.300 ;
        RECT 1413.180 2.890 1420.980 4.300 ;
        RECT 1422.140 2.890 1429.940 4.300 ;
        RECT 1431.100 2.890 1438.900 4.300 ;
        RECT 1440.060 2.890 1447.860 4.300 ;
        RECT 1449.020 2.890 1456.820 4.300 ;
        RECT 1457.980 2.890 1465.780 4.300 ;
        RECT 1466.940 2.890 1474.740 4.300 ;
        RECT 1475.900 2.890 1483.700 4.300 ;
        RECT 1484.860 2.890 1492.660 4.300 ;
        RECT 1493.820 2.890 1501.620 4.300 ;
        RECT 1502.780 2.890 1510.580 4.300 ;
        RECT 1511.740 2.890 1519.540 4.300 ;
        RECT 1520.700 2.890 1528.500 4.300 ;
        RECT 1529.660 2.890 1537.460 4.300 ;
        RECT 1538.620 2.890 1546.420 4.300 ;
        RECT 1547.580 2.890 1555.380 4.300 ;
        RECT 1556.540 2.890 1564.340 4.300 ;
        RECT 1565.500 2.890 1573.300 4.300 ;
        RECT 1574.460 2.890 1582.260 4.300 ;
        RECT 1583.420 2.890 1591.220 4.300 ;
        RECT 1592.380 2.890 1600.180 4.300 ;
        RECT 1601.340 2.890 1609.140 4.300 ;
        RECT 1610.300 2.890 1618.100 4.300 ;
        RECT 1619.260 2.890 1627.060 4.300 ;
        RECT 1628.220 2.890 1636.020 4.300 ;
        RECT 1637.180 2.890 1644.980 4.300 ;
        RECT 1646.140 2.890 1653.940 4.300 ;
        RECT 1655.100 2.890 1662.900 4.300 ;
        RECT 1664.060 2.890 1671.860 4.300 ;
        RECT 1673.020 2.890 1680.820 4.300 ;
        RECT 1681.980 2.890 1689.780 4.300 ;
        RECT 1690.940 2.890 1698.740 4.300 ;
        RECT 1699.900 2.890 1707.700 4.300 ;
        RECT 1708.860 2.890 1716.660 4.300 ;
        RECT 1717.820 2.890 1725.620 4.300 ;
        RECT 1726.780 2.890 1734.580 4.300 ;
        RECT 1735.740 2.890 1743.540 4.300 ;
        RECT 1744.700 2.890 1752.500 4.300 ;
        RECT 1753.660 2.890 1761.460 4.300 ;
        RECT 1762.620 2.890 1770.420 4.300 ;
        RECT 1771.580 2.890 1779.380 4.300 ;
        RECT 1780.540 2.890 1788.340 4.300 ;
        RECT 1789.500 2.890 1797.300 4.300 ;
        RECT 1798.460 2.890 1806.260 4.300 ;
        RECT 1807.420 2.890 1815.220 4.300 ;
        RECT 1816.380 2.890 1824.180 4.300 ;
        RECT 1825.340 2.890 1833.140 4.300 ;
        RECT 1834.300 2.890 1842.100 4.300 ;
        RECT 1843.260 2.890 1851.060 4.300 ;
        RECT 1852.220 2.890 1860.020 4.300 ;
        RECT 1861.180 2.890 1868.980 4.300 ;
        RECT 1870.140 2.890 1877.940 4.300 ;
        RECT 1879.100 2.890 1886.900 4.300 ;
        RECT 1888.060 2.890 1895.860 4.300 ;
        RECT 1897.020 2.890 1904.820 4.300 ;
        RECT 1905.980 2.890 1913.780 4.300 ;
        RECT 1914.940 2.890 1922.740 4.300 ;
        RECT 1923.900 2.890 1931.700 4.300 ;
        RECT 1932.860 2.890 1940.660 4.300 ;
        RECT 1941.820 2.890 1949.620 4.300 ;
        RECT 1950.780 2.890 1958.580 4.300 ;
        RECT 1959.740 2.890 1967.540 4.300 ;
        RECT 1968.700 2.890 1976.500 4.300 ;
        RECT 1977.660 2.890 1985.460 4.300 ;
        RECT 1986.620 2.890 1994.420 4.300 ;
        RECT 1995.580 2.890 2003.380 4.300 ;
        RECT 2004.540 2.890 2012.340 4.300 ;
        RECT 2013.500 2.890 2021.300 4.300 ;
        RECT 2022.460 2.890 2030.260 4.300 ;
        RECT 2031.420 2.890 2039.220 4.300 ;
        RECT 2040.380 2.890 2048.180 4.300 ;
        RECT 2049.340 2.890 2057.140 4.300 ;
        RECT 2058.300 2.890 2066.100 4.300 ;
        RECT 2067.260 2.890 2075.060 4.300 ;
        RECT 2076.220 2.890 2084.020 4.300 ;
        RECT 2085.180 2.890 2092.980 4.300 ;
        RECT 2094.140 2.890 2101.940 4.300 ;
        RECT 2103.100 2.890 2110.900 4.300 ;
        RECT 2112.060 2.890 2119.860 4.300 ;
        RECT 2121.020 2.890 2128.820 4.300 ;
        RECT 2129.980 2.890 2137.780 4.300 ;
        RECT 2138.940 2.890 2146.740 4.300 ;
        RECT 2147.900 2.890 2155.700 4.300 ;
        RECT 2156.860 2.890 2164.660 4.300 ;
        RECT 2165.820 2.890 2173.620 4.300 ;
        RECT 2174.780 2.890 2182.580 4.300 ;
        RECT 2183.740 2.890 2191.540 4.300 ;
        RECT 2192.700 2.890 2200.500 4.300 ;
        RECT 2201.660 2.890 2209.460 4.300 ;
        RECT 2210.620 2.890 2218.420 4.300 ;
        RECT 2219.580 2.890 2227.380 4.300 ;
        RECT 2228.540 2.890 2236.340 4.300 ;
        RECT 2237.500 2.890 2245.300 4.300 ;
        RECT 2246.460 2.890 2254.260 4.300 ;
        RECT 2255.420 2.890 2263.220 4.300 ;
        RECT 2264.380 2.890 2272.180 4.300 ;
        RECT 2273.340 2.890 2281.140 4.300 ;
        RECT 2282.300 2.890 2290.100 4.300 ;
        RECT 2291.260 2.890 2299.060 4.300 ;
        RECT 2300.220 2.890 2308.020 4.300 ;
        RECT 2309.180 2.890 2316.980 4.300 ;
        RECT 2318.140 2.890 2325.940 4.300 ;
        RECT 2327.100 2.890 2334.900 4.300 ;
        RECT 2336.060 2.890 2343.860 4.300 ;
        RECT 2345.020 2.890 2352.820 4.300 ;
        RECT 2353.980 2.890 2361.780 4.300 ;
        RECT 2362.940 2.890 2370.740 4.300 ;
        RECT 2371.900 2.890 2379.700 4.300 ;
        RECT 2380.860 2.890 2388.660 4.300 ;
        RECT 2389.820 2.890 2397.620 4.300 ;
        RECT 2398.780 2.890 2406.580 4.300 ;
        RECT 2407.740 2.890 2415.540 4.300 ;
        RECT 2416.700 2.890 2424.500 4.300 ;
        RECT 2425.660 2.890 2433.460 4.300 ;
        RECT 2434.620 2.890 2442.420 4.300 ;
        RECT 2443.580 2.890 2451.380 4.300 ;
        RECT 2452.540 2.890 2460.340 4.300 ;
        RECT 2461.500 2.890 2469.300 4.300 ;
        RECT 2470.460 2.890 2478.260 4.300 ;
        RECT 2479.420 2.890 2487.220 4.300 ;
        RECT 2488.380 2.890 2496.180 4.300 ;
        RECT 2497.340 2.890 2505.140 4.300 ;
        RECT 2506.300 2.890 2514.100 4.300 ;
        RECT 2515.260 2.890 2523.060 4.300 ;
        RECT 2524.220 2.890 2532.020 4.300 ;
        RECT 2533.180 2.890 2540.980 4.300 ;
        RECT 2542.140 2.890 2549.940 4.300 ;
        RECT 2551.100 2.890 2558.900 4.300 ;
        RECT 2560.060 2.890 2567.860 4.300 ;
        RECT 2569.020 2.890 2576.820 4.300 ;
        RECT 2577.980 2.890 2585.780 4.300 ;
        RECT 2586.940 2.890 2594.740 4.300 ;
        RECT 2595.900 2.890 2603.700 4.300 ;
        RECT 2604.860 2.890 2612.660 4.300 ;
        RECT 2613.820 2.890 2621.620 4.300 ;
        RECT 2622.780 2.890 2630.580 4.300 ;
        RECT 2631.740 2.890 2639.540 4.300 ;
        RECT 2640.700 2.890 2648.500 4.300 ;
        RECT 2649.660 2.890 2657.460 4.300 ;
        RECT 2658.620 2.890 2666.420 4.300 ;
        RECT 2667.580 2.890 2675.380 4.300 ;
        RECT 2676.540 2.890 2684.340 4.300 ;
        RECT 2685.500 2.890 2693.300 4.300 ;
        RECT 2694.460 2.890 2702.260 4.300 ;
        RECT 2703.420 2.890 2711.220 4.300 ;
        RECT 2712.380 2.890 2720.180 4.300 ;
        RECT 2721.340 2.890 2729.140 4.300 ;
        RECT 2730.300 2.890 2738.100 4.300 ;
        RECT 2739.260 2.890 2747.060 4.300 ;
        RECT 2748.220 2.890 2756.020 4.300 ;
        RECT 2757.180 2.890 2764.980 4.300 ;
        RECT 2766.140 2.890 2773.940 4.300 ;
        RECT 2775.100 2.890 2782.900 4.300 ;
        RECT 2784.060 2.890 2863.700 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 2842.300 2866.470 2874.340 ;
        RECT 4.000 2841.140 2866.170 2842.300 ;
        RECT 4.000 2838.940 2866.470 2841.140 ;
        RECT 4.300 2837.780 2866.470 2838.940 ;
        RECT 4.000 2788.540 2866.470 2837.780 ;
        RECT 4.000 2787.380 2866.170 2788.540 ;
        RECT 4.000 2786.300 2866.470 2787.380 ;
        RECT 4.300 2785.140 2866.470 2786.300 ;
        RECT 4.000 2734.780 2866.470 2785.140 ;
        RECT 4.000 2733.660 2866.170 2734.780 ;
        RECT 4.300 2733.620 2866.170 2733.660 ;
        RECT 4.300 2732.500 2866.470 2733.620 ;
        RECT 4.000 2681.020 2866.470 2732.500 ;
        RECT 4.300 2679.860 2866.170 2681.020 ;
        RECT 4.000 2628.380 2866.470 2679.860 ;
        RECT 4.300 2627.260 2866.470 2628.380 ;
        RECT 4.300 2627.220 2866.170 2627.260 ;
        RECT 4.000 2626.100 2866.170 2627.220 ;
        RECT 4.000 2575.740 2866.470 2626.100 ;
        RECT 4.300 2574.580 2866.470 2575.740 ;
        RECT 4.000 2573.500 2866.470 2574.580 ;
        RECT 4.000 2572.340 2866.170 2573.500 ;
        RECT 4.000 2523.100 2866.470 2572.340 ;
        RECT 4.300 2521.940 2866.470 2523.100 ;
        RECT 4.000 2519.740 2866.470 2521.940 ;
        RECT 4.000 2518.580 2866.170 2519.740 ;
        RECT 4.000 2470.460 2866.470 2518.580 ;
        RECT 4.300 2469.300 2866.470 2470.460 ;
        RECT 4.000 2465.980 2866.470 2469.300 ;
        RECT 4.000 2464.820 2866.170 2465.980 ;
        RECT 4.000 2417.820 2866.470 2464.820 ;
        RECT 4.300 2416.660 2866.470 2417.820 ;
        RECT 4.000 2412.220 2866.470 2416.660 ;
        RECT 4.000 2411.060 2866.170 2412.220 ;
        RECT 4.000 2365.180 2866.470 2411.060 ;
        RECT 4.300 2364.020 2866.470 2365.180 ;
        RECT 4.000 2358.460 2866.470 2364.020 ;
        RECT 4.000 2357.300 2866.170 2358.460 ;
        RECT 4.000 2312.540 2866.470 2357.300 ;
        RECT 4.300 2311.380 2866.470 2312.540 ;
        RECT 4.000 2304.700 2866.470 2311.380 ;
        RECT 4.000 2303.540 2866.170 2304.700 ;
        RECT 4.000 2259.900 2866.470 2303.540 ;
        RECT 4.300 2258.740 2866.470 2259.900 ;
        RECT 4.000 2250.940 2866.470 2258.740 ;
        RECT 4.000 2249.780 2866.170 2250.940 ;
        RECT 4.000 2207.260 2866.470 2249.780 ;
        RECT 4.300 2206.100 2866.470 2207.260 ;
        RECT 4.000 2197.180 2866.470 2206.100 ;
        RECT 4.000 2196.020 2866.170 2197.180 ;
        RECT 4.000 2154.620 2866.470 2196.020 ;
        RECT 4.300 2153.460 2866.470 2154.620 ;
        RECT 4.000 2143.420 2866.470 2153.460 ;
        RECT 4.000 2142.260 2866.170 2143.420 ;
        RECT 4.000 2101.980 2866.470 2142.260 ;
        RECT 4.300 2100.820 2866.470 2101.980 ;
        RECT 4.000 2089.660 2866.470 2100.820 ;
        RECT 4.000 2088.500 2866.170 2089.660 ;
        RECT 4.000 2049.340 2866.470 2088.500 ;
        RECT 4.300 2048.180 2866.470 2049.340 ;
        RECT 4.000 2035.900 2866.470 2048.180 ;
        RECT 4.000 2034.740 2866.170 2035.900 ;
        RECT 4.000 1996.700 2866.470 2034.740 ;
        RECT 4.300 1995.540 2866.470 1996.700 ;
        RECT 4.000 1982.140 2866.470 1995.540 ;
        RECT 4.000 1980.980 2866.170 1982.140 ;
        RECT 4.000 1944.060 2866.470 1980.980 ;
        RECT 4.300 1942.900 2866.470 1944.060 ;
        RECT 4.000 1928.380 2866.470 1942.900 ;
        RECT 4.000 1927.220 2866.170 1928.380 ;
        RECT 4.000 1891.420 2866.470 1927.220 ;
        RECT 4.300 1890.260 2866.470 1891.420 ;
        RECT 4.000 1874.620 2866.470 1890.260 ;
        RECT 4.000 1873.460 2866.170 1874.620 ;
        RECT 4.000 1838.780 2866.470 1873.460 ;
        RECT 4.300 1837.620 2866.470 1838.780 ;
        RECT 4.000 1820.860 2866.470 1837.620 ;
        RECT 4.000 1819.700 2866.170 1820.860 ;
        RECT 4.000 1786.140 2866.470 1819.700 ;
        RECT 4.300 1784.980 2866.470 1786.140 ;
        RECT 4.000 1767.100 2866.470 1784.980 ;
        RECT 4.000 1765.940 2866.170 1767.100 ;
        RECT 4.000 1733.500 2866.470 1765.940 ;
        RECT 4.300 1732.340 2866.470 1733.500 ;
        RECT 4.000 1713.340 2866.470 1732.340 ;
        RECT 4.000 1712.180 2866.170 1713.340 ;
        RECT 4.000 1680.860 2866.470 1712.180 ;
        RECT 4.300 1679.700 2866.470 1680.860 ;
        RECT 4.000 1659.580 2866.470 1679.700 ;
        RECT 4.000 1658.420 2866.170 1659.580 ;
        RECT 4.000 1628.220 2866.470 1658.420 ;
        RECT 4.300 1627.060 2866.470 1628.220 ;
        RECT 4.000 1605.820 2866.470 1627.060 ;
        RECT 4.000 1604.660 2866.170 1605.820 ;
        RECT 4.000 1575.580 2866.470 1604.660 ;
        RECT 4.300 1574.420 2866.470 1575.580 ;
        RECT 4.000 1552.060 2866.470 1574.420 ;
        RECT 4.000 1550.900 2866.170 1552.060 ;
        RECT 4.000 1522.940 2866.470 1550.900 ;
        RECT 4.300 1521.780 2866.470 1522.940 ;
        RECT 4.000 1498.300 2866.470 1521.780 ;
        RECT 4.000 1497.140 2866.170 1498.300 ;
        RECT 4.000 1470.300 2866.470 1497.140 ;
        RECT 4.300 1469.140 2866.470 1470.300 ;
        RECT 4.000 1444.540 2866.470 1469.140 ;
        RECT 4.000 1443.380 2866.170 1444.540 ;
        RECT 4.000 1417.660 2866.470 1443.380 ;
        RECT 4.300 1416.500 2866.470 1417.660 ;
        RECT 4.000 1390.780 2866.470 1416.500 ;
        RECT 4.000 1389.620 2866.170 1390.780 ;
        RECT 4.000 1365.020 2866.470 1389.620 ;
        RECT 4.300 1363.860 2866.470 1365.020 ;
        RECT 4.000 1337.020 2866.470 1363.860 ;
        RECT 4.000 1335.860 2866.170 1337.020 ;
        RECT 4.000 1312.380 2866.470 1335.860 ;
        RECT 4.300 1311.220 2866.470 1312.380 ;
        RECT 4.000 1283.260 2866.470 1311.220 ;
        RECT 4.000 1282.100 2866.170 1283.260 ;
        RECT 4.000 1259.740 2866.470 1282.100 ;
        RECT 4.300 1258.580 2866.470 1259.740 ;
        RECT 4.000 1229.500 2866.470 1258.580 ;
        RECT 4.000 1228.340 2866.170 1229.500 ;
        RECT 4.000 1207.100 2866.470 1228.340 ;
        RECT 4.300 1205.940 2866.470 1207.100 ;
        RECT 4.000 1175.740 2866.470 1205.940 ;
        RECT 4.000 1174.580 2866.170 1175.740 ;
        RECT 4.000 1154.460 2866.470 1174.580 ;
        RECT 4.300 1153.300 2866.470 1154.460 ;
        RECT 4.000 1121.980 2866.470 1153.300 ;
        RECT 4.000 1120.820 2866.170 1121.980 ;
        RECT 4.000 1101.820 2866.470 1120.820 ;
        RECT 4.300 1100.660 2866.470 1101.820 ;
        RECT 4.000 1068.220 2866.470 1100.660 ;
        RECT 4.000 1067.060 2866.170 1068.220 ;
        RECT 4.000 1049.180 2866.470 1067.060 ;
        RECT 4.300 1048.020 2866.470 1049.180 ;
        RECT 4.000 1014.460 2866.470 1048.020 ;
        RECT 4.000 1013.300 2866.170 1014.460 ;
        RECT 4.000 996.540 2866.470 1013.300 ;
        RECT 4.300 995.380 2866.470 996.540 ;
        RECT 4.000 960.700 2866.470 995.380 ;
        RECT 4.000 959.540 2866.170 960.700 ;
        RECT 4.000 943.900 2866.470 959.540 ;
        RECT 4.300 942.740 2866.470 943.900 ;
        RECT 4.000 906.940 2866.470 942.740 ;
        RECT 4.000 905.780 2866.170 906.940 ;
        RECT 4.000 891.260 2866.470 905.780 ;
        RECT 4.300 890.100 2866.470 891.260 ;
        RECT 4.000 853.180 2866.470 890.100 ;
        RECT 4.000 852.020 2866.170 853.180 ;
        RECT 4.000 838.620 2866.470 852.020 ;
        RECT 4.300 837.460 2866.470 838.620 ;
        RECT 4.000 799.420 2866.470 837.460 ;
        RECT 4.000 798.260 2866.170 799.420 ;
        RECT 4.000 785.980 2866.470 798.260 ;
        RECT 4.300 784.820 2866.470 785.980 ;
        RECT 4.000 745.660 2866.470 784.820 ;
        RECT 4.000 744.500 2866.170 745.660 ;
        RECT 4.000 733.340 2866.470 744.500 ;
        RECT 4.300 732.180 2866.470 733.340 ;
        RECT 4.000 691.900 2866.470 732.180 ;
        RECT 4.000 690.740 2866.170 691.900 ;
        RECT 4.000 680.700 2866.470 690.740 ;
        RECT 4.300 679.540 2866.470 680.700 ;
        RECT 4.000 638.140 2866.470 679.540 ;
        RECT 4.000 636.980 2866.170 638.140 ;
        RECT 4.000 628.060 2866.470 636.980 ;
        RECT 4.300 626.900 2866.470 628.060 ;
        RECT 4.000 584.380 2866.470 626.900 ;
        RECT 4.000 583.220 2866.170 584.380 ;
        RECT 4.000 575.420 2866.470 583.220 ;
        RECT 4.300 574.260 2866.470 575.420 ;
        RECT 4.000 530.620 2866.470 574.260 ;
        RECT 4.000 529.460 2866.170 530.620 ;
        RECT 4.000 522.780 2866.470 529.460 ;
        RECT 4.300 521.620 2866.470 522.780 ;
        RECT 4.000 476.860 2866.470 521.620 ;
        RECT 4.000 475.700 2866.170 476.860 ;
        RECT 4.000 470.140 2866.470 475.700 ;
        RECT 4.300 468.980 2866.470 470.140 ;
        RECT 4.000 423.100 2866.470 468.980 ;
        RECT 4.000 421.940 2866.170 423.100 ;
        RECT 4.000 417.500 2866.470 421.940 ;
        RECT 4.300 416.340 2866.470 417.500 ;
        RECT 4.000 369.340 2866.470 416.340 ;
        RECT 4.000 368.180 2866.170 369.340 ;
        RECT 4.000 364.860 2866.470 368.180 ;
        RECT 4.300 363.700 2866.470 364.860 ;
        RECT 4.000 315.580 2866.470 363.700 ;
        RECT 4.000 314.420 2866.170 315.580 ;
        RECT 4.000 312.220 2866.470 314.420 ;
        RECT 4.300 311.060 2866.470 312.220 ;
        RECT 4.000 261.820 2866.470 311.060 ;
        RECT 4.000 260.660 2866.170 261.820 ;
        RECT 4.000 259.580 2866.470 260.660 ;
        RECT 4.300 258.420 2866.470 259.580 ;
        RECT 4.000 208.060 2866.470 258.420 ;
        RECT 4.000 206.940 2866.170 208.060 ;
        RECT 4.300 206.900 2866.170 206.940 ;
        RECT 4.300 205.780 2866.470 206.900 ;
        RECT 4.000 154.300 2866.470 205.780 ;
        RECT 4.300 153.140 2866.170 154.300 ;
        RECT 4.000 101.660 2866.470 153.140 ;
        RECT 4.300 100.540 2866.470 101.660 ;
        RECT 4.300 100.500 2866.170 100.540 ;
        RECT 4.000 99.380 2866.170 100.500 ;
        RECT 4.000 49.020 2866.470 99.380 ;
        RECT 4.300 47.860 2866.470 49.020 ;
        RECT 4.000 46.780 2866.470 47.860 ;
        RECT 4.000 45.620 2866.170 46.780 ;
        RECT 4.000 2.940 2866.470 45.620 ;
      LAYER Metal4 ;
        RECT 10.220 2870.040 2855.860 2874.390 ;
        RECT 10.220 15.080 21.940 2870.040 ;
        RECT 24.140 15.080 98.740 2870.040 ;
        RECT 100.940 15.080 175.540 2870.040 ;
        RECT 177.740 15.080 252.340 2870.040 ;
        RECT 254.540 15.080 329.140 2870.040 ;
        RECT 331.340 15.080 405.940 2870.040 ;
        RECT 408.140 15.080 482.740 2870.040 ;
        RECT 484.940 15.080 559.540 2870.040 ;
        RECT 561.740 15.080 636.340 2870.040 ;
        RECT 638.540 15.080 713.140 2870.040 ;
        RECT 715.340 15.080 789.940 2870.040 ;
        RECT 792.140 15.080 866.740 2870.040 ;
        RECT 868.940 15.080 943.540 2870.040 ;
        RECT 945.740 15.080 1020.340 2870.040 ;
        RECT 1022.540 15.080 1097.140 2870.040 ;
        RECT 1099.340 15.080 1173.940 2870.040 ;
        RECT 1176.140 15.080 1250.740 2870.040 ;
        RECT 1252.940 15.080 1327.540 2870.040 ;
        RECT 1329.740 15.080 1404.340 2870.040 ;
        RECT 1406.540 15.080 1481.140 2870.040 ;
        RECT 1483.340 15.080 1557.940 2870.040 ;
        RECT 1560.140 15.080 1634.740 2870.040 ;
        RECT 1636.940 15.080 1711.540 2870.040 ;
        RECT 1713.740 15.080 1788.340 2870.040 ;
        RECT 1790.540 15.080 1865.140 2870.040 ;
        RECT 1867.340 15.080 1941.940 2870.040 ;
        RECT 1944.140 15.080 2018.740 2870.040 ;
        RECT 2020.940 15.080 2095.540 2870.040 ;
        RECT 2097.740 15.080 2172.340 2870.040 ;
        RECT 2174.540 15.080 2249.140 2870.040 ;
        RECT 2251.340 15.080 2325.940 2870.040 ;
        RECT 2328.140 15.080 2402.740 2870.040 ;
        RECT 2404.940 15.080 2479.540 2870.040 ;
        RECT 2481.740 15.080 2556.340 2870.040 ;
        RECT 2558.540 15.080 2633.140 2870.040 ;
        RECT 2635.340 15.080 2709.940 2870.040 ;
        RECT 2712.140 15.080 2786.740 2870.040 ;
        RECT 2788.940 15.080 2855.860 2870.040 ;
        RECT 10.220 6.810 2855.860 15.080 ;
  END
END rift2Wrap
END LIBRARY

