magic
tech gf180mcuD
magscale 1 10
timestamp 1698902861
<< metal2 >>
rect 11032 595672 11256 597000
rect 11032 595560 11284 595672
rect 11228 588868 11284 595560
rect 32396 595644 33012 595700
rect 33096 595672 33320 597000
rect 55160 595672 55384 597000
rect 11228 588802 11284 588812
rect 16492 588868 16548 588878
rect 16492 585592 16548 588812
rect 32396 585592 32452 595644
rect 32956 595476 33012 595644
rect 33068 595560 33320 595672
rect 55132 595560 55384 595672
rect 77224 595672 77448 597000
rect 99288 595672 99512 597000
rect 121352 595672 121576 597000
rect 77224 595560 77476 595672
rect 33068 595476 33124 595560
rect 32956 595420 33124 595476
rect 48300 591332 48356 591342
rect 48300 585592 48356 591276
rect 55132 591332 55188 595560
rect 55132 591266 55188 591276
rect 77420 591332 77476 595560
rect 99260 595560 99512 595672
rect 121324 595560 121576 595672
rect 143416 595672 143640 597000
rect 165480 595672 165704 597000
rect 187544 595672 187768 597000
rect 209608 595672 209832 597000
rect 231672 595672 231896 597000
rect 253736 595672 253960 597000
rect 275800 595672 276024 597000
rect 297864 595672 298088 597000
rect 319928 595672 320152 597000
rect 341992 595672 342216 597000
rect 364056 595672 364280 597000
rect 386120 595672 386344 597000
rect 143416 595560 143668 595672
rect 77420 591266 77476 591276
rect 80108 591332 80164 591342
rect 80108 585592 80164 591276
rect 96012 591332 96068 591342
rect 96012 585592 96068 591276
rect 99260 591332 99316 595560
rect 99260 591266 99316 591276
rect 111916 588868 111972 588878
rect 111916 585592 111972 588812
rect 121324 588868 121380 595560
rect 121324 588802 121380 588812
rect 143612 588028 143668 595560
rect 165452 595560 165704 595672
rect 187516 595560 187768 595672
rect 209580 595560 209832 595672
rect 231644 595560 231896 595672
rect 253708 595560 253960 595672
rect 275772 595560 276024 595672
rect 297836 595560 298088 595672
rect 319900 595560 320152 595672
rect 341964 595560 342216 595672
rect 364028 595560 364280 595672
rect 386092 595560 386344 595672
rect 408184 595560 408408 597000
rect 430248 595672 430472 597000
rect 452312 595672 452536 597000
rect 474376 595672 474600 597000
rect 496440 595672 496664 597000
rect 518504 595672 518728 597000
rect 540568 595672 540792 597000
rect 562632 595672 562856 597000
rect 584696 595672 584920 597000
rect 430220 595560 430472 595672
rect 452284 595560 452536 595672
rect 474348 595560 474600 595672
rect 496412 595560 496664 595672
rect 518476 595560 518728 595672
rect 540540 595560 540792 595672
rect 562604 595560 562856 595672
rect 584668 595560 584920 595672
rect 159628 590548 159684 590558
rect 143612 587972 143780 588028
rect 143724 585592 143780 587972
rect 159628 585592 159684 590492
rect 165452 590548 165508 595560
rect 165452 590482 165508 590492
rect 175532 588868 175588 588878
rect 175532 585592 175588 588812
rect 187516 588868 187572 595560
rect 187516 588802 187572 588812
rect 207340 591332 207396 591342
rect 207340 585592 207396 591276
rect 209580 591332 209636 595560
rect 209580 591266 209636 591276
rect 223244 590548 223300 590558
rect 223244 585592 223300 590492
rect 231644 590548 231700 595560
rect 231644 590482 231700 590492
rect 239148 588868 239204 588878
rect 239148 585592 239204 588812
rect 253708 588868 253764 595560
rect 253708 588802 253764 588812
rect 270956 591332 271012 591342
rect 270956 585592 271012 591276
rect 275772 591332 275828 595560
rect 275772 591266 275828 591276
rect 286860 588868 286916 588878
rect 286860 585592 286916 588812
rect 297836 588868 297892 595560
rect 297836 588802 297892 588812
rect 302764 588868 302820 588878
rect 302764 585592 302820 588812
rect 319900 588868 319956 595560
rect 319900 588802 319956 588812
rect 334572 590548 334628 590558
rect 334572 585592 334628 590492
rect 341964 590548 342020 595560
rect 341964 590482 342020 590492
rect 350476 590548 350532 590558
rect 350476 585592 350532 590492
rect 364028 590548 364084 595560
rect 364028 590482 364084 590492
rect 366380 588868 366436 588878
rect 366380 585592 366436 588812
rect 386092 588868 386148 595560
rect 386092 588802 386148 588812
rect 398188 588868 398244 588878
rect 398188 585592 398244 588812
rect 408268 588868 408324 595560
rect 429996 590548 430052 590558
rect 408268 588802 408324 588812
rect 414092 588868 414148 588878
rect 414092 585592 414148 588812
rect 429996 585592 430052 590492
rect 430220 588868 430276 595560
rect 452284 590548 452340 595560
rect 452284 590482 452340 590492
rect 461804 590548 461860 590558
rect 430220 588802 430276 588812
rect 461804 585592 461860 590492
rect 474348 590548 474404 595560
rect 474348 590482 474404 590492
rect 493612 590548 493668 590558
rect 477708 588868 477764 588878
rect 477708 585592 477764 588812
rect 493612 585592 493668 590492
rect 496412 588868 496468 595560
rect 518476 590548 518532 595560
rect 518476 590482 518532 590492
rect 496412 588802 496468 588812
rect 525420 588868 525476 588878
rect 525420 585592 525476 588812
rect 540540 588868 540596 595560
rect 540540 588802 540596 588812
rect 541324 590660 541380 590670
rect 541324 585592 541380 590604
rect 562604 590660 562660 595560
rect 562604 590594 562660 590604
rect 557228 590548 557284 590558
rect 557228 585592 557284 590492
rect 584668 590548 584724 595560
rect 584668 590482 584724 590492
rect 11564 5908 11620 5918
rect 11564 480 11620 5852
rect 25228 5908 25284 8120
rect 25228 5842 25284 5852
rect 26796 5012 26852 5022
rect 24892 4900 24948 4910
rect 22988 4788 23044 4798
rect 21084 4676 21140 4686
rect 19180 4564 19236 4574
rect 17276 4452 17332 4462
rect 15372 4340 15428 4350
rect 13356 4228 13412 4238
rect 13356 480 13412 4172
rect 15372 480 15428 4284
rect 17276 480 17332 4396
rect 19180 480 19236 4508
rect 21084 480 21140 4620
rect 22988 480 23044 4732
rect 24892 480 24948 4844
rect 26796 480 26852 4956
rect 27020 4228 27076 8120
rect 28812 4340 28868 8120
rect 30604 4452 30660 8120
rect 32396 4564 32452 8120
rect 34188 4676 34244 8120
rect 35980 4788 36036 8120
rect 37772 4900 37828 8120
rect 39564 5012 39620 8120
rect 39564 4946 39620 4956
rect 37772 4834 37828 4844
rect 35980 4722 36036 4732
rect 40124 4788 40180 4798
rect 34188 4610 34244 4620
rect 38220 4676 38276 4686
rect 32396 4498 32452 4508
rect 36316 4564 36372 4574
rect 30604 4386 30660 4396
rect 34412 4452 34468 4462
rect 28812 4274 28868 4284
rect 32508 4340 32564 4350
rect 27020 4162 27076 4172
rect 30604 4228 30660 4238
rect 28700 4116 28756 4126
rect 28700 480 28756 4060
rect 30604 480 30660 4172
rect 32508 480 32564 4284
rect 34412 480 34468 4396
rect 36316 480 36372 4508
rect 38220 480 38276 4620
rect 40124 480 40180 4732
rect 41356 4116 41412 8120
rect 41356 4050 41412 4060
rect 41916 4900 41972 4910
rect 41916 480 41972 4844
rect 43148 4228 43204 8120
rect 44940 4340 44996 8120
rect 46732 4452 46788 8120
rect 48524 4564 48580 8120
rect 50316 4676 50372 8120
rect 52108 4788 52164 8120
rect 53900 4900 53956 8120
rect 53900 4834 53956 4844
rect 55356 4900 55412 4910
rect 52108 4722 52164 4732
rect 53452 4788 53508 4798
rect 50316 4610 50372 4620
rect 51548 4676 51604 4686
rect 48524 4498 48580 4508
rect 49644 4564 49700 4574
rect 46732 4386 46788 4396
rect 47740 4452 47796 4462
rect 44940 4274 44996 4284
rect 45836 4340 45892 4350
rect 43148 4162 43204 4172
rect 43932 4228 43988 4238
rect 43932 480 43988 4172
rect 45836 480 45892 4284
rect 47740 480 47796 4396
rect 49644 480 49700 4508
rect 51548 480 51604 4620
rect 53452 480 53508 4732
rect 55356 480 55412 4844
rect 55692 4228 55748 8120
rect 57484 4340 57540 8120
rect 59276 4452 59332 8120
rect 61068 4564 61124 8120
rect 62860 4676 62916 8120
rect 64652 4788 64708 8120
rect 64652 4722 64708 4732
rect 64876 5012 64932 5022
rect 62860 4610 62916 4620
rect 61068 4498 61124 4508
rect 62972 4564 63028 4574
rect 59276 4386 59332 4396
rect 61180 4452 61236 4462
rect 57484 4274 57540 4284
rect 55692 4162 55748 4172
rect 57260 4228 57316 4238
rect 57260 480 57316 4172
rect 59164 4116 59220 4126
rect 59164 480 59220 4060
rect 61180 2212 61236 4396
rect 61068 2156 61236 2212
rect 61068 480 61124 2156
rect 62972 480 63028 4508
rect 64876 480 64932 4956
rect 66444 4900 66500 8120
rect 66444 4834 66500 4844
rect 66780 4676 66836 4686
rect 66780 480 66836 4620
rect 68236 4228 68292 8120
rect 68236 4162 68292 4172
rect 68684 4228 68740 4238
rect 68684 480 68740 4172
rect 70028 4116 70084 8120
rect 71820 4452 71876 8120
rect 73612 4564 73668 8120
rect 75404 5012 75460 8120
rect 75404 4946 75460 4956
rect 76300 4788 76356 4798
rect 73612 4498 73668 4508
rect 74396 4564 74452 4574
rect 71820 4386 71876 4396
rect 72492 4452 72548 4462
rect 70028 4050 70084 4060
rect 70476 4340 70532 4350
rect 70476 480 70532 4284
rect 72492 480 72548 4396
rect 74396 480 74452 4508
rect 76300 480 76356 4732
rect 77196 4676 77252 8120
rect 77196 4610 77252 4620
rect 78204 4676 78260 4686
rect 78204 480 78260 4620
rect 78988 4228 79044 8120
rect 80780 4340 80836 8120
rect 82572 4452 82628 8120
rect 84364 4564 84420 8120
rect 86156 4788 86212 8120
rect 86156 4722 86212 4732
rect 87724 4788 87780 4798
rect 84364 4498 84420 4508
rect 85820 4564 85876 4574
rect 82572 4386 82628 4396
rect 80780 4274 80836 4284
rect 82012 4340 82068 4350
rect 78988 4162 79044 4172
rect 80108 4228 80164 4238
rect 80108 480 80164 4172
rect 82012 480 82068 4284
rect 83916 4116 83972 4126
rect 83916 480 83972 4060
rect 85820 480 85876 4508
rect 87724 480 87780 4732
rect 87948 4676 88004 8120
rect 87948 4610 88004 4620
rect 89628 4676 89684 4686
rect 89628 480 89684 4620
rect 89740 4228 89796 8120
rect 90860 8092 91560 8148
rect 90860 4340 90916 8092
rect 90860 4274 90916 4284
rect 89740 4162 89796 4172
rect 91532 4228 91588 4238
rect 91532 480 91588 4172
rect 93324 4116 93380 8120
rect 95116 4564 95172 8120
rect 96908 4788 96964 8120
rect 96908 4722 96964 4732
rect 98700 4676 98756 8120
rect 98700 4610 98756 4620
rect 95116 4498 95172 4508
rect 99036 4564 99092 4574
rect 97244 4452 97300 4462
rect 93324 4050 93380 4060
rect 93436 4340 93492 4350
rect 93436 480 93492 4284
rect 95340 4116 95396 4126
rect 95340 480 95396 4060
rect 97244 480 97300 4396
rect 99036 480 99092 4508
rect 100492 4228 100548 8120
rect 102284 4340 102340 8120
rect 102284 4274 102340 4284
rect 102956 4340 103012 4350
rect 100492 4162 100548 4172
rect 101052 4228 101108 4238
rect 101052 480 101108 4172
rect 102956 480 103012 4284
rect 104076 4116 104132 8120
rect 104076 4050 104132 4060
rect 104860 4676 104916 4686
rect 104860 480 104916 4620
rect 105868 4452 105924 8120
rect 107660 4564 107716 8120
rect 107660 4498 107716 4508
rect 105868 4386 105924 4396
rect 109452 4228 109508 8120
rect 111244 4340 111300 8120
rect 113036 4676 113092 8120
rect 113036 4610 113092 4620
rect 114380 4676 114436 4686
rect 111244 4274 111300 4284
rect 112476 4340 112532 4350
rect 109452 4162 109508 4172
rect 110572 4228 110628 4238
rect 108668 4116 108724 4126
rect 106764 4004 106820 4014
rect 106764 480 106820 3948
rect 108668 480 108724 4060
rect 110572 480 110628 4172
rect 112476 480 112532 4284
rect 114380 480 114436 4620
rect 114828 4004 114884 8120
rect 114828 3938 114884 3948
rect 116284 4452 116340 4462
rect 116284 480 116340 4396
rect 116620 4116 116676 8120
rect 118412 4228 118468 8120
rect 120204 4340 120260 8120
rect 121996 4676 122052 8120
rect 121996 4610 122052 4620
rect 123788 4452 123844 8120
rect 123788 4386 123844 4396
rect 123900 4676 123956 4686
rect 120204 4274 120260 4284
rect 118412 4162 118468 4172
rect 116620 4050 116676 4060
rect 121996 4116 122052 4126
rect 120092 4004 120148 4014
rect 118188 3892 118244 3902
rect 118188 480 118244 3836
rect 120092 480 120148 3948
rect 121996 480 122052 4060
rect 123900 480 123956 4620
rect 125580 3892 125636 8120
rect 125580 3826 125636 3836
rect 125804 4788 125860 4798
rect 125804 480 125860 4732
rect 127372 4004 127428 8120
rect 127372 3938 127428 3948
rect 127596 4452 127652 4462
rect 127596 480 127652 4396
rect 129164 4116 129220 8120
rect 130956 4676 131012 8120
rect 132748 4788 132804 8120
rect 132748 4722 132804 4732
rect 130956 4610 131012 4620
rect 134540 4452 134596 8120
rect 134540 4386 134596 4396
rect 135324 4452 135380 4462
rect 129164 4050 129220 4060
rect 129612 4228 129668 4238
rect 129612 480 129668 4172
rect 133420 4116 133476 4126
rect 131516 4004 131572 4014
rect 131516 480 131572 3948
rect 133420 480 133476 4060
rect 135324 480 135380 4396
rect 136332 4228 136388 8120
rect 136332 4162 136388 4172
rect 137228 4228 137284 4238
rect 137228 480 137284 4172
rect 138124 4004 138180 8120
rect 138124 3938 138180 3948
rect 139132 4340 139188 4350
rect 139132 480 139188 4284
rect 139916 4116 139972 8120
rect 139916 4050 139972 4060
rect 141036 4564 141092 4574
rect 141036 480 141092 4508
rect 141708 4452 141764 8120
rect 141708 4386 141764 4396
rect 143500 4228 143556 8120
rect 145292 4340 145348 8120
rect 145292 4274 145348 4284
rect 146748 4676 146804 4686
rect 143500 4162 143556 4172
rect 144844 4116 144900 4126
rect 142940 4004 142996 4014
rect 142940 480 142996 3948
rect 144844 480 144900 4060
rect 146748 480 146804 4620
rect 147084 4564 147140 8120
rect 147084 4498 147140 4508
rect 148652 4564 148708 4574
rect 148652 480 148708 4508
rect 148876 4004 148932 8120
rect 148876 3938 148932 3948
rect 150556 4452 150612 4462
rect 150556 480 150612 4396
rect 150668 4116 150724 8120
rect 152460 4676 152516 8120
rect 152460 4610 152516 4620
rect 154252 4564 154308 8120
rect 154252 4498 154308 4508
rect 156044 4452 156100 8120
rect 156044 4386 156100 4396
rect 150668 4050 150724 4060
rect 152460 4228 152516 4238
rect 152460 480 152516 4172
rect 157836 4228 157892 8120
rect 157836 4162 157892 4172
rect 158172 4116 158228 4126
rect 156156 4004 156212 4014
rect 154364 3892 154420 3902
rect 154364 480 154420 3836
rect 156156 480 156212 3948
rect 158172 480 158228 4060
rect 159628 3892 159684 8120
rect 159628 3826 159684 3836
rect 160076 4228 160132 4238
rect 160076 480 160132 4172
rect 161420 4004 161476 8120
rect 161420 3938 161476 3948
rect 161980 4340 162036 4350
rect 161980 480 162036 4284
rect 163212 4116 163268 8120
rect 163212 4050 163268 4060
rect 163884 4452 163940 4462
rect 163884 480 163940 4396
rect 165004 4228 165060 8120
rect 166796 4340 166852 8120
rect 168588 4452 168644 8120
rect 168588 4386 168644 4396
rect 166796 4274 166852 4284
rect 165004 4162 165060 4172
rect 165788 4228 165844 4238
rect 165788 480 165844 4172
rect 170380 4228 170436 8120
rect 170380 4162 170436 4172
rect 171500 5124 171556 5134
rect 169596 4116 169652 4126
rect 167692 4004 167748 4014
rect 167692 480 167748 3948
rect 169596 480 169652 4060
rect 171500 480 171556 5068
rect 172172 4004 172228 8120
rect 172172 3938 172228 3948
rect 173404 6020 173460 6030
rect 173404 480 173460 5964
rect 173964 4116 174020 8120
rect 173964 4050 174020 4060
rect 175308 6132 175364 6142
rect 175308 480 175364 6076
rect 175756 5124 175812 8120
rect 177548 6020 177604 8120
rect 179340 6132 179396 8120
rect 179340 6066 179396 6076
rect 177548 5954 177604 5964
rect 175756 5058 175812 5068
rect 177212 5348 177268 5358
rect 177212 480 177268 5292
rect 181132 5348 181188 8120
rect 181132 5282 181188 5292
rect 179116 5236 179172 5246
rect 179116 480 179172 5180
rect 182924 5236 182980 8120
rect 182924 5170 182980 5180
rect 181020 5124 181076 5134
rect 181020 480 181076 5068
rect 184716 5124 184772 8120
rect 184716 5058 184772 5068
rect 184716 4340 184772 4350
rect 182924 4116 182980 4126
rect 182924 480 182980 4060
rect 184716 480 184772 4284
rect 186508 4116 186564 8120
rect 186508 4050 186564 4060
rect 186732 5908 186788 5918
rect 186732 480 186788 5852
rect 188300 4340 188356 8120
rect 190092 5908 190148 8120
rect 190092 5842 190148 5852
rect 190540 5236 190596 5246
rect 188300 4274 188356 4284
rect 188636 5124 188692 5134
rect 188636 480 188692 5068
rect 190540 480 190596 5180
rect 191884 5124 191940 8120
rect 193676 5236 193732 8120
rect 193676 5170 193732 5180
rect 194348 5236 194404 5246
rect 191884 5058 191940 5068
rect 192444 5124 192500 5134
rect 192444 480 192500 5068
rect 194348 480 194404 5180
rect 195468 5124 195524 8120
rect 197260 5236 197316 8120
rect 197260 5170 197316 5180
rect 198156 5908 198212 5918
rect 195468 5058 195524 5068
rect 196252 5124 196308 5134
rect 196252 480 196308 5068
rect 198156 480 198212 5852
rect 199052 5124 199108 8120
rect 200844 5908 200900 8120
rect 200844 5842 200900 5852
rect 199052 5058 199108 5068
rect 200060 5236 200116 5246
rect 200060 480 200116 5180
rect 202636 5236 202692 8120
rect 202636 5170 202692 5180
rect 203868 5236 203924 5246
rect 201964 5124 202020 5134
rect 201964 480 202020 5068
rect 203868 480 203924 5180
rect 204428 5124 204484 8120
rect 206220 5236 206276 8120
rect 206220 5170 206276 5180
rect 207676 5236 207732 5246
rect 204428 5058 204484 5068
rect 205772 5124 205828 5134
rect 205772 480 205828 5068
rect 207676 480 207732 5180
rect 208012 5124 208068 8120
rect 209804 5236 209860 8120
rect 209804 5170 209860 5180
rect 211484 6020 211540 6030
rect 208012 5058 208068 5068
rect 209580 5124 209636 5134
rect 209580 480 209636 5068
rect 211484 480 211540 5964
rect 211596 5124 211652 8120
rect 213388 6020 213444 8120
rect 213388 5954 213444 5964
rect 211596 5058 211652 5068
rect 213276 5236 213332 5246
rect 213276 480 213332 5180
rect 215180 5236 215236 8120
rect 215180 5170 215236 5180
rect 215292 5124 215348 5134
rect 215292 480 215348 5068
rect 216972 5124 217028 8120
rect 216972 5058 217028 5068
rect 217196 5124 217252 5134
rect 217196 480 217252 5068
rect 218764 5124 218820 8120
rect 220108 8092 220584 8148
rect 221788 8092 222376 8148
rect 220108 5124 220164 8092
rect 221788 5124 221844 8092
rect 218764 5058 218820 5068
rect 219884 5068 220164 5124
rect 221676 5068 221844 5124
rect 222908 5908 222964 5918
rect 219100 480 219268 532
rect 11368 392 11620 480
rect 11368 -960 11592 392
rect 13272 -960 13496 480
rect 15176 392 15428 480
rect 17080 392 17332 480
rect 18984 392 19236 480
rect 20888 392 21140 480
rect 22792 392 23044 480
rect 24696 392 24948 480
rect 26600 392 26852 480
rect 28504 392 28756 480
rect 30408 392 30660 480
rect 32312 392 32564 480
rect 34216 392 34468 480
rect 36120 392 36372 480
rect 38024 392 38276 480
rect 39928 392 40180 480
rect 15176 -960 15400 392
rect 17080 -960 17304 392
rect 18984 -960 19208 392
rect 20888 -960 21112 392
rect 22792 -960 23016 392
rect 24696 -960 24920 392
rect 26600 -960 26824 392
rect 28504 -960 28728 392
rect 30408 -960 30632 392
rect 32312 -960 32536 392
rect 34216 -960 34440 392
rect 36120 -960 36344 392
rect 38024 -960 38248 392
rect 39928 -960 40152 392
rect 41832 -960 42056 480
rect 43736 392 43988 480
rect 45640 392 45892 480
rect 47544 392 47796 480
rect 49448 392 49700 480
rect 51352 392 51604 480
rect 53256 392 53508 480
rect 55160 392 55412 480
rect 57064 392 57316 480
rect 58968 392 59220 480
rect 60872 392 61124 480
rect 62776 392 63028 480
rect 64680 392 64932 480
rect 66584 392 66836 480
rect 68488 392 68740 480
rect 43736 -960 43960 392
rect 45640 -960 45864 392
rect 47544 -960 47768 392
rect 49448 -960 49672 392
rect 51352 -960 51576 392
rect 53256 -960 53480 392
rect 55160 -960 55384 392
rect 57064 -960 57288 392
rect 58968 -960 59192 392
rect 60872 -960 61096 392
rect 62776 -960 63000 392
rect 64680 -960 64904 392
rect 66584 -960 66808 392
rect 68488 -960 68712 392
rect 70392 -960 70616 480
rect 72296 392 72548 480
rect 74200 392 74452 480
rect 76104 392 76356 480
rect 78008 392 78260 480
rect 79912 392 80164 480
rect 81816 392 82068 480
rect 83720 392 83972 480
rect 85624 392 85876 480
rect 87528 392 87780 480
rect 89432 392 89684 480
rect 91336 392 91588 480
rect 93240 392 93492 480
rect 95144 392 95396 480
rect 97048 392 97300 480
rect 72296 -960 72520 392
rect 74200 -960 74424 392
rect 76104 -960 76328 392
rect 78008 -960 78232 392
rect 79912 -960 80136 392
rect 81816 -960 82040 392
rect 83720 -960 83944 392
rect 85624 -960 85848 392
rect 87528 -960 87752 392
rect 89432 -960 89656 392
rect 91336 -960 91560 392
rect 93240 -960 93464 392
rect 95144 -960 95368 392
rect 97048 -960 97272 392
rect 98952 -960 99176 480
rect 100856 392 101108 480
rect 102760 392 103012 480
rect 104664 392 104916 480
rect 106568 392 106820 480
rect 108472 392 108724 480
rect 110376 392 110628 480
rect 112280 392 112532 480
rect 114184 392 114436 480
rect 116088 392 116340 480
rect 117992 392 118244 480
rect 119896 392 120148 480
rect 121800 392 122052 480
rect 123704 392 123956 480
rect 125608 392 125860 480
rect 100856 -960 101080 392
rect 102760 -960 102984 392
rect 104664 -960 104888 392
rect 106568 -960 106792 392
rect 108472 -960 108696 392
rect 110376 -960 110600 392
rect 112280 -960 112504 392
rect 114184 -960 114408 392
rect 116088 -960 116312 392
rect 117992 -960 118216 392
rect 119896 -960 120120 392
rect 121800 -960 122024 392
rect 123704 -960 123928 392
rect 125608 -960 125832 392
rect 127512 -960 127736 480
rect 129416 392 129668 480
rect 131320 392 131572 480
rect 133224 392 133476 480
rect 135128 392 135380 480
rect 137032 392 137284 480
rect 138936 392 139188 480
rect 140840 392 141092 480
rect 142744 392 142996 480
rect 144648 392 144900 480
rect 146552 392 146804 480
rect 148456 392 148708 480
rect 150360 392 150612 480
rect 152264 392 152516 480
rect 154168 392 154420 480
rect 129416 -960 129640 392
rect 131320 -960 131544 392
rect 133224 -960 133448 392
rect 135128 -960 135352 392
rect 137032 -960 137256 392
rect 138936 -960 139160 392
rect 140840 -960 141064 392
rect 142744 -960 142968 392
rect 144648 -960 144872 392
rect 146552 -960 146776 392
rect 148456 -960 148680 392
rect 150360 -960 150584 392
rect 152264 -960 152488 392
rect 154168 -960 154392 392
rect 156072 -960 156296 480
rect 157976 392 158228 480
rect 159880 392 160132 480
rect 161784 392 162036 480
rect 163688 392 163940 480
rect 165592 392 165844 480
rect 167496 392 167748 480
rect 169400 392 169652 480
rect 171304 392 171556 480
rect 173208 392 173460 480
rect 175112 392 175364 480
rect 177016 392 177268 480
rect 178920 392 179172 480
rect 180824 392 181076 480
rect 182728 392 182980 480
rect 157976 -960 158200 392
rect 159880 -960 160104 392
rect 161784 -960 162008 392
rect 163688 -960 163912 392
rect 165592 -960 165816 392
rect 167496 -960 167720 392
rect 169400 -960 169624 392
rect 171304 -960 171528 392
rect 173208 -960 173432 392
rect 175112 -960 175336 392
rect 177016 -960 177240 392
rect 178920 -960 179144 392
rect 180824 -960 181048 392
rect 182728 -960 182952 392
rect 184632 -960 184856 480
rect 186536 392 186788 480
rect 188440 392 188692 480
rect 190344 392 190596 480
rect 192248 392 192500 480
rect 194152 392 194404 480
rect 196056 392 196308 480
rect 197960 392 198212 480
rect 199864 392 200116 480
rect 201768 392 202020 480
rect 203672 392 203924 480
rect 205576 392 205828 480
rect 207480 392 207732 480
rect 209384 392 209636 480
rect 211288 392 211540 480
rect 186536 -960 186760 392
rect 188440 -960 188664 392
rect 190344 -960 190568 392
rect 192248 -960 192472 392
rect 194152 -960 194376 392
rect 196056 -960 196280 392
rect 197960 -960 198184 392
rect 199864 -960 200088 392
rect 201768 -960 201992 392
rect 203672 -960 203896 392
rect 205576 -960 205800 392
rect 207480 -960 207704 392
rect 209384 -960 209608 392
rect 211288 -960 211512 392
rect 213192 -960 213416 480
rect 215096 392 215348 480
rect 217000 392 217252 480
rect 218904 476 219268 480
rect 218904 392 219156 476
rect 219212 420 219268 476
rect 219884 420 219940 5068
rect 221004 480 221172 532
rect 215096 -960 215320 392
rect 217000 -960 217224 392
rect 218904 -960 219128 392
rect 219212 364 219940 420
rect 220808 476 221172 480
rect 220808 392 221060 476
rect 221116 420 221172 476
rect 221676 420 221732 5068
rect 222908 480 222964 5852
rect 224140 5908 224196 8120
rect 224140 5842 224196 5852
rect 225148 8092 225960 8148
rect 226828 8092 227752 8148
rect 228620 8092 229544 8148
rect 230524 8092 231336 8148
rect 232428 8092 233128 8148
rect 234332 8092 234920 8148
rect 236236 8092 236712 8148
rect 238140 8092 238504 8148
rect 225148 5124 225204 8092
rect 226828 5124 226884 8092
rect 224812 5068 225204 5124
rect 226716 5068 226884 5124
rect 224812 480 224868 5068
rect 226716 480 226772 5068
rect 228620 480 228676 8092
rect 230524 480 230580 8092
rect 232428 480 232484 8092
rect 234332 480 234388 8092
rect 236236 480 236292 8092
rect 238140 480 238196 8092
rect 240268 5124 240324 8120
rect 241948 8092 242088 8148
rect 241948 5124 242004 8092
rect 240044 5068 240324 5124
rect 241836 5068 242004 5124
rect 240044 480 240100 5068
rect 241836 480 241892 5068
rect 243852 480 243908 8120
rect 245644 480 245700 8120
rect 247436 480 247492 8120
rect 249256 8092 249396 8148
rect 251048 8092 251300 8148
rect 252840 8092 253204 8148
rect 254632 8092 255108 8148
rect 256424 8092 257012 8148
rect 249340 480 249396 8092
rect 251244 480 251300 8092
rect 253148 480 253204 8092
rect 255052 480 255108 8092
rect 256956 5124 257012 8092
rect 258188 5908 258244 8120
rect 260008 8092 260372 8148
rect 261800 8092 262052 8148
rect 263592 8092 263732 8148
rect 258188 5842 258244 5852
rect 258860 5908 258916 5918
rect 256956 5068 257124 5124
rect 257068 480 257124 5068
rect 258860 480 258916 5852
rect 260316 5124 260372 8092
rect 261996 5124 262052 8092
rect 263676 5124 263732 8092
rect 265356 5124 265412 8120
rect 267176 8092 267876 8148
rect 268968 8092 269668 8148
rect 260316 5068 260484 5124
rect 261996 5068 262164 5124
rect 263676 5068 263844 5124
rect 220808 -960 221032 392
rect 221116 364 221732 420
rect 222712 392 222964 480
rect 224616 392 224868 480
rect 226520 392 226772 480
rect 228424 392 228676 480
rect 230328 392 230580 480
rect 232232 392 232484 480
rect 234136 392 234388 480
rect 236040 392 236292 480
rect 237944 392 238196 480
rect 239848 392 240100 480
rect 222712 -960 222936 392
rect 224616 -960 224840 392
rect 226520 -960 226744 392
rect 228424 -960 228648 392
rect 230328 -960 230552 392
rect 232232 -960 232456 392
rect 234136 -960 234360 392
rect 236040 -960 236264 392
rect 237944 -960 238168 392
rect 239848 -960 240072 392
rect 241752 -960 241976 480
rect 243656 392 243908 480
rect 243656 -960 243880 392
rect 245560 -960 245784 480
rect 247436 392 247688 480
rect 249340 392 249592 480
rect 251244 392 251496 480
rect 253148 392 253400 480
rect 255052 392 255304 480
rect 247464 -960 247688 392
rect 249368 -960 249592 392
rect 251272 -960 251496 392
rect 253176 -960 253400 392
rect 255080 -960 255304 392
rect 256984 -960 257208 480
rect 258860 392 259112 480
rect 258888 -960 259112 392
rect 260428 420 260484 5068
rect 260652 480 260820 532
rect 260652 476 261016 480
rect 260652 420 260708 476
rect 260428 364 260708 420
rect 260764 392 261016 476
rect 260792 -960 261016 392
rect 262108 420 262164 5068
rect 262556 480 262724 532
rect 262556 476 262920 480
rect 262556 420 262612 476
rect 262108 364 262612 420
rect 262668 392 262920 476
rect 262696 -960 262920 392
rect 263788 420 263844 5068
rect 265356 5058 265412 5068
rect 266476 5124 266532 5134
rect 264460 480 264628 532
rect 266476 480 266532 5068
rect 264460 476 264824 480
rect 264460 420 264516 476
rect 263788 364 264516 420
rect 264572 392 264824 476
rect 266476 392 266728 480
rect 264600 -960 264824 392
rect 266504 -960 266728 392
rect 267820 420 267876 8092
rect 268268 480 268436 532
rect 268268 476 268632 480
rect 268268 420 268324 476
rect 267820 364 268324 420
rect 268380 392 268632 476
rect 268408 -960 268632 392
rect 269612 420 269668 8092
rect 270732 5124 270788 8120
rect 270732 5058 270788 5068
rect 272188 5124 272244 5134
rect 270172 480 270340 532
rect 272188 480 272244 5068
rect 272524 5124 272580 8120
rect 272524 5058 272580 5068
rect 274092 5124 274148 5134
rect 274092 480 274148 5068
rect 274316 5124 274372 8120
rect 276108 5236 276164 8120
rect 277900 5460 277956 8120
rect 277900 5394 277956 5404
rect 276108 5170 276164 5180
rect 277900 5236 277956 5246
rect 274316 5058 274372 5068
rect 275996 5124 276052 5134
rect 275996 480 276052 5068
rect 277900 480 277956 5180
rect 279692 5124 279748 8120
rect 281484 5908 281540 8120
rect 281484 5842 281540 5852
rect 279692 5058 279748 5068
rect 279804 5460 279860 5470
rect 279804 480 279860 5404
rect 281708 5124 281764 5134
rect 281708 480 281764 5068
rect 283276 4116 283332 8120
rect 283276 4050 283332 4060
rect 283612 5908 283668 5918
rect 283612 480 283668 5852
rect 285068 4004 285124 8120
rect 285068 3938 285124 3948
rect 285628 4116 285684 4126
rect 285628 480 285684 4060
rect 286860 4116 286916 8120
rect 286860 4050 286916 4060
rect 287420 4004 287476 4014
rect 287420 480 287476 3948
rect 288652 4004 288708 8120
rect 288652 3938 288708 3948
rect 289324 4116 289380 4126
rect 289324 480 289380 4060
rect 290444 4116 290500 8120
rect 292236 4228 292292 8120
rect 294028 5124 294084 8120
rect 295820 5236 295876 8120
rect 295820 5170 295876 5180
rect 294028 5058 294084 5068
rect 296940 5124 296996 5134
rect 292236 4162 292292 4172
rect 295036 4228 295092 4238
rect 290444 4050 290500 4060
rect 293132 4116 293188 4126
rect 291228 4004 291284 4014
rect 291228 480 291284 3948
rect 293132 480 293188 4060
rect 295036 480 295092 4172
rect 296940 480 296996 5068
rect 297612 4116 297668 8120
rect 297612 4050 297668 4060
rect 298844 5236 298900 5246
rect 298844 480 298900 5180
rect 299404 4004 299460 8120
rect 299404 3938 299460 3948
rect 300748 4116 300804 4126
rect 300748 480 300804 4060
rect 301196 4116 301252 8120
rect 302988 4228 303044 8120
rect 304780 4452 304836 8120
rect 304780 4386 304836 4396
rect 302988 4162 303044 4172
rect 306460 4228 306516 4238
rect 301196 4050 301252 4060
rect 304556 4116 304612 4126
rect 302652 4004 302708 4014
rect 302652 480 302708 3948
rect 304556 480 304612 4060
rect 306460 480 306516 4172
rect 306572 4116 306628 8120
rect 308364 4676 308420 8120
rect 310156 5124 310212 8120
rect 311948 5236 312004 8120
rect 313740 5908 313796 8120
rect 315532 6132 315588 8120
rect 315532 6066 315588 6076
rect 317324 6020 317380 8120
rect 317324 5954 317380 5964
rect 313740 5842 313796 5852
rect 317884 5908 317940 5918
rect 311948 5170 312004 5180
rect 315980 5236 316036 5246
rect 310156 5058 310212 5068
rect 314188 5124 314244 5134
rect 308364 4610 308420 4620
rect 312172 4676 312228 4686
rect 306572 4050 306628 4060
rect 308364 4452 308420 4462
rect 308364 480 308420 4396
rect 310268 4116 310324 4126
rect 310268 480 310324 4060
rect 312172 480 312228 4620
rect 314188 480 314244 5068
rect 315980 480 316036 5180
rect 317884 480 317940 5852
rect 319116 5124 319172 8120
rect 319116 5058 319172 5068
rect 319788 6132 319844 6142
rect 319788 480 319844 6076
rect 320908 4116 320964 8120
rect 320908 4050 320964 4060
rect 321692 6020 321748 6030
rect 321692 480 321748 5964
rect 322700 4004 322756 8120
rect 324492 6020 324548 8120
rect 324492 5954 324548 5964
rect 326284 5908 326340 8120
rect 328076 6132 328132 8120
rect 328076 6066 328132 6076
rect 326284 5842 326340 5852
rect 329308 6020 329364 6030
rect 322700 3938 322756 3948
rect 323596 5124 323652 5134
rect 323596 480 323652 5068
rect 325500 4116 325556 4126
rect 325500 480 325556 4060
rect 327404 4004 327460 4014
rect 327404 480 327460 3948
rect 329308 480 329364 5964
rect 329868 5124 329924 8120
rect 329868 5058 329924 5068
rect 331212 5908 331268 5918
rect 331212 480 331268 5852
rect 331660 5236 331716 8120
rect 331660 5170 331716 5180
rect 333116 6132 333172 6142
rect 333116 480 333172 6076
rect 333452 5348 333508 8120
rect 333452 5282 333508 5292
rect 335020 5124 335076 5134
rect 335020 480 335076 5068
rect 335244 5124 335300 8120
rect 337036 6132 337092 8120
rect 337036 6066 337092 6076
rect 338828 6020 338884 8120
rect 338828 5954 338884 5964
rect 340620 5908 340676 8120
rect 340620 5842 340676 5852
rect 338828 5348 338884 5358
rect 335244 5058 335300 5068
rect 336924 5236 336980 5246
rect 336924 480 336980 5180
rect 338828 480 338884 5292
rect 340732 5124 340788 5134
rect 340732 480 340788 5068
rect 342412 5124 342468 8120
rect 342412 5058 342468 5068
rect 342748 6132 342804 6142
rect 342748 480 342804 6076
rect 344204 5236 344260 8120
rect 344204 5170 344260 5180
rect 344540 6020 344596 6030
rect 344540 480 344596 5964
rect 345996 5348 346052 8120
rect 345996 5282 346052 5292
rect 346444 5908 346500 5918
rect 346444 480 346500 5852
rect 347788 5908 347844 8120
rect 349580 6244 349636 8120
rect 349580 6178 349636 6188
rect 351372 6132 351428 8120
rect 351372 6066 351428 6076
rect 347788 5842 347844 5852
rect 352156 5348 352212 5358
rect 350252 5236 350308 5246
rect 348348 5124 348404 5134
rect 348348 480 348404 5068
rect 350252 480 350308 5180
rect 352156 480 352212 5292
rect 353164 5124 353220 8120
rect 353164 5058 353220 5068
rect 354060 5908 354116 5918
rect 354060 480 354116 5852
rect 354956 5236 355012 8120
rect 354956 5170 355012 5180
rect 355964 6244 356020 6254
rect 355964 480 356020 6188
rect 356748 5348 356804 8120
rect 356748 5282 356804 5292
rect 357868 6132 357924 6142
rect 357868 480 357924 6076
rect 358540 6132 358596 8120
rect 358540 6066 358596 6076
rect 360332 6020 360388 8120
rect 360332 5954 360388 5964
rect 362124 5908 362180 8120
rect 362124 5842 362180 5852
rect 363580 5348 363636 5358
rect 361676 5236 361732 5246
rect 359772 5124 359828 5134
rect 359772 480 359828 5068
rect 361676 480 361732 5180
rect 363580 480 363636 5292
rect 363916 4452 363972 8120
rect 363916 4386 363972 4396
rect 365484 6132 365540 6142
rect 365484 480 365540 6076
rect 365708 4116 365764 8120
rect 365708 4050 365764 4060
rect 367388 6020 367444 6030
rect 367388 480 367444 5964
rect 367500 4004 367556 8120
rect 369320 8092 369572 8148
rect 367500 3938 367556 3948
rect 369292 5908 369348 5918
rect 369292 480 369348 5852
rect 369516 4340 369572 8092
rect 369516 4274 369572 4284
rect 371084 4228 371140 8120
rect 371084 4162 371140 4172
rect 371308 4452 371364 4462
rect 371308 480 371364 4396
rect 372876 4452 372932 8120
rect 374668 6020 374724 8120
rect 374668 5954 374724 5964
rect 376460 5124 376516 8120
rect 376460 5058 376516 5068
rect 372876 4386 372932 4396
rect 376908 4340 376964 4350
rect 373100 4116 373156 4126
rect 373100 480 373156 4060
rect 375004 4004 375060 4014
rect 375004 480 375060 3948
rect 376908 480 376964 4284
rect 378252 4116 378308 8120
rect 378252 4050 378308 4060
rect 378812 4228 378868 4238
rect 378812 480 378868 4172
rect 380044 4228 380100 8120
rect 381836 4676 381892 8120
rect 381836 4610 381892 4620
rect 382620 6020 382676 6030
rect 380044 4162 380100 4172
rect 380716 4452 380772 4462
rect 380716 480 380772 4396
rect 382620 480 382676 5964
rect 383628 4564 383684 8120
rect 383628 4498 383684 4508
rect 384524 5124 384580 5134
rect 384524 480 384580 5068
rect 385420 4452 385476 8120
rect 385420 4386 385476 4396
rect 387212 4340 387268 8120
rect 387212 4274 387268 4284
rect 388332 4228 388388 4238
rect 386428 4116 386484 4126
rect 386428 480 386484 4060
rect 388332 480 388388 4172
rect 389004 4116 389060 8120
rect 390796 6356 390852 8120
rect 392588 6468 392644 8120
rect 392588 6402 392644 6412
rect 390796 6290 390852 6300
rect 394380 5908 394436 8120
rect 396172 6244 396228 8120
rect 396172 6178 396228 6188
rect 397964 6132 398020 8120
rect 397964 6066 398020 6076
rect 399756 6020 399812 8120
rect 399756 5954 399812 5964
rect 399868 6356 399924 6366
rect 394380 5842 394436 5852
rect 389004 4050 389060 4060
rect 390236 4676 390292 4686
rect 390236 480 390292 4620
rect 392140 4564 392196 4574
rect 392140 480 392196 4508
rect 394044 4452 394100 4462
rect 394044 480 394100 4396
rect 395948 4340 396004 4350
rect 395948 480 396004 4284
rect 397852 4116 397908 4126
rect 397852 480 397908 4060
rect 399868 480 399924 6300
rect 401548 4116 401604 8120
rect 401548 4050 401604 4060
rect 401660 6468 401716 6478
rect 401660 480 401716 6412
rect 403340 4228 403396 8120
rect 403340 4162 403396 4172
rect 403564 5908 403620 5918
rect 403564 480 403620 5852
rect 405132 5908 405188 8120
rect 406924 6356 406980 8120
rect 408716 6468 408772 8120
rect 408716 6402 408772 6412
rect 406924 6290 406980 6300
rect 405132 5842 405188 5852
rect 405468 6244 405524 6254
rect 405468 480 405524 6188
rect 410508 6244 410564 8120
rect 410508 6178 410564 6188
rect 407372 6132 407428 6142
rect 407372 480 407428 6076
rect 409276 6020 409332 6030
rect 409276 480 409332 5964
rect 412300 5124 412356 8120
rect 414092 6020 414148 8120
rect 414092 5954 414148 5964
rect 412300 5058 412356 5068
rect 414988 5908 415044 5918
rect 413084 4228 413140 4238
rect 411180 4116 411236 4126
rect 411180 480 411236 4060
rect 413084 480 413140 4172
rect 414988 480 415044 5852
rect 415884 5908 415940 8120
rect 415884 5842 415940 5852
rect 416892 6356 416948 6366
rect 416892 480 416948 6300
rect 417676 6356 417732 8120
rect 419468 6692 419524 8120
rect 419468 6626 419524 6636
rect 417676 6290 417732 6300
rect 418796 6468 418852 6478
rect 418796 480 418852 6412
rect 421260 6468 421316 8120
rect 423052 6580 423108 8120
rect 423052 6514 423108 6524
rect 421260 6402 421316 6412
rect 420700 6244 420756 6254
rect 420700 480 420756 6188
rect 424844 6244 424900 8120
rect 424844 6178 424900 6188
rect 426636 6132 426692 8120
rect 428456 8092 429156 8148
rect 426636 6066 426692 6076
rect 428428 6356 428484 6366
rect 424508 6020 424564 6030
rect 422604 5124 422660 5134
rect 422604 480 422660 5068
rect 424508 480 424564 5964
rect 426412 5908 426468 5918
rect 426412 480 426468 5852
rect 428428 480 428484 6300
rect 429100 6020 429156 8092
rect 429100 5954 429156 5964
rect 430220 5908 430276 8120
rect 430220 5842 430276 5852
rect 430332 6692 430388 6702
rect 430332 480 430388 6636
rect 432012 6356 432068 8120
rect 432012 6290 432068 6300
rect 432124 6468 432180 6478
rect 432124 480 432180 6412
rect 433804 6468 433860 8120
rect 433804 6402 433860 6412
rect 434028 6580 434084 6590
rect 434028 480 434084 6524
rect 435596 6580 435652 8120
rect 435596 6514 435652 6524
rect 435932 6244 435988 6254
rect 435932 480 435988 6188
rect 437388 6244 437444 8120
rect 437388 6178 437444 6188
rect 437836 6132 437892 6142
rect 437836 480 437892 6076
rect 439180 6132 439236 8120
rect 439180 6066 439236 6076
rect 439740 6020 439796 6030
rect 439740 480 439796 5964
rect 440972 6020 441028 8120
rect 440972 5954 441028 5964
rect 441644 5908 441700 5918
rect 441644 480 441700 5852
rect 442764 5908 442820 8120
rect 442764 5842 442820 5852
rect 443548 6356 443604 6366
rect 443548 480 443604 6300
rect 444556 6356 444612 8120
rect 444556 6290 444612 6300
rect 445452 6468 445508 6478
rect 445452 480 445508 6412
rect 446348 6468 446404 8120
rect 446348 6402 446404 6412
rect 447356 6580 447412 6590
rect 447356 480 447412 6524
rect 448140 5796 448196 8120
rect 448140 5730 448196 5740
rect 449260 6244 449316 6254
rect 449260 480 449316 6188
rect 449932 6244 449988 8120
rect 449932 6178 449988 6188
rect 451164 6132 451220 6142
rect 451164 480 451220 6076
rect 451724 6132 451780 8120
rect 451724 6066 451780 6076
rect 453068 6020 453124 6030
rect 453068 480 453124 5964
rect 453516 6020 453572 8120
rect 453516 5954 453572 5964
rect 454972 5908 455028 5918
rect 454972 480 455028 5852
rect 455308 5908 455364 8120
rect 457100 6692 457156 8120
rect 457100 6626 457156 6636
rect 458892 6580 458948 8120
rect 458892 6514 458948 6524
rect 458780 6468 458836 6478
rect 455308 5842 455364 5852
rect 456988 6356 457044 6366
rect 456988 480 457044 6300
rect 458780 480 458836 6412
rect 460684 6468 460740 8120
rect 460684 6402 460740 6412
rect 462476 6356 462532 8120
rect 462476 6290 462532 6300
rect 462588 6244 462644 6254
rect 460684 5796 460740 5806
rect 460684 480 460740 5740
rect 462588 480 462644 6188
rect 464268 6244 464324 8120
rect 464268 6178 464324 6188
rect 464492 6132 464548 6142
rect 464492 480 464548 6076
rect 466060 6132 466116 8120
rect 466060 6066 466116 6076
rect 466396 6020 466452 6030
rect 466396 480 466452 5964
rect 467852 6020 467908 8120
rect 467852 5954 467908 5964
rect 468300 5908 468356 5918
rect 468300 480 468356 5852
rect 469644 5908 469700 8120
rect 469644 5842 469700 5852
rect 470204 6692 470260 6702
rect 470204 480 470260 6636
rect 471436 4676 471492 8120
rect 471436 4610 471492 4620
rect 472108 6580 472164 6590
rect 472108 480 472164 6524
rect 473228 4788 473284 8120
rect 473228 4722 473284 4732
rect 474012 6468 474068 6478
rect 474012 480 474068 6412
rect 475020 4564 475076 8120
rect 475020 4498 475076 4508
rect 475916 6356 475972 6366
rect 475916 480 475972 6300
rect 476812 4340 476868 8120
rect 476812 4274 476868 4284
rect 477820 6244 477876 6254
rect 477820 480 477876 6188
rect 478604 4228 478660 8120
rect 478604 4162 478660 4172
rect 479724 6132 479780 6142
rect 479724 480 479780 6076
rect 480396 4452 480452 8120
rect 480396 4386 480452 4396
rect 481628 6020 481684 6030
rect 481628 480 481684 5964
rect 482188 6020 482244 8120
rect 482188 5954 482244 5964
rect 483532 5908 483588 5918
rect 483532 480 483588 5852
rect 483980 5908 484036 8120
rect 483980 5842 484036 5852
rect 485772 4900 485828 8120
rect 485772 4834 485828 4844
rect 487340 4788 487396 4798
rect 485548 4676 485604 4686
rect 485548 480 485604 4620
rect 487340 480 487396 4732
rect 487564 4788 487620 8120
rect 487564 4722 487620 4732
rect 489356 4676 489412 8120
rect 489356 4610 489412 4620
rect 489244 4564 489300 4574
rect 489244 480 489300 4508
rect 491148 4564 491204 8120
rect 491148 4498 491204 4508
rect 491148 4340 491204 4350
rect 491148 480 491204 4284
rect 492940 4340 492996 8120
rect 492940 4274 492996 4284
rect 493052 4228 493108 4238
rect 493052 480 493108 4172
rect 494732 4228 494788 8120
rect 494732 4162 494788 4172
rect 494956 4452 495012 4462
rect 494956 480 495012 4396
rect 496524 4452 496580 8120
rect 498316 6356 498372 8120
rect 500108 6468 500164 8120
rect 500108 6402 500164 6412
rect 498316 6290 498372 6300
rect 501900 6244 501956 8120
rect 501900 6178 501956 6188
rect 503692 6132 503748 8120
rect 503692 6066 503748 6076
rect 496524 4386 496580 4396
rect 496860 6020 496916 6030
rect 496860 480 496916 5964
rect 505484 6020 505540 8120
rect 505484 5954 505540 5964
rect 498764 5908 498820 5918
rect 498764 480 498820 5852
rect 507276 5908 507332 8120
rect 507276 5842 507332 5852
rect 500668 4900 500724 4910
rect 500668 480 500724 4844
rect 502572 4788 502628 4798
rect 502572 480 502628 4732
rect 504476 4676 504532 4686
rect 504476 480 504532 4620
rect 506380 4564 506436 4574
rect 506380 480 506436 4508
rect 508284 4340 508340 4350
rect 508284 480 508340 4284
rect 509068 4340 509124 8120
rect 509068 4274 509124 4284
rect 510188 4228 510244 4238
rect 510188 480 510244 4172
rect 510860 4228 510916 8120
rect 512652 5796 512708 8120
rect 514444 6580 514500 8120
rect 516236 6692 516292 8120
rect 516236 6626 516292 6636
rect 514444 6514 514500 6524
rect 515900 6468 515956 6478
rect 512652 5730 512708 5740
rect 514108 6356 514164 6366
rect 510860 4162 510916 4172
rect 512092 4452 512148 4462
rect 512092 480 512148 4396
rect 514108 480 514164 6300
rect 515900 480 515956 6412
rect 518028 6468 518084 8120
rect 518028 6402 518084 6412
rect 519820 6356 519876 8120
rect 519820 6290 519876 6300
rect 517804 6244 517860 6254
rect 517804 480 517860 6188
rect 521612 6244 521668 8120
rect 521612 6178 521668 6188
rect 519708 6132 519764 6142
rect 519708 480 519764 6076
rect 523404 6132 523460 8120
rect 523404 6066 523460 6076
rect 521612 6020 521668 6030
rect 521612 480 521668 5964
rect 523516 5908 523572 5918
rect 523516 480 523572 5852
rect 525196 4676 525252 8120
rect 526988 6020 527044 8120
rect 526988 5954 527044 5964
rect 528780 5908 528836 8120
rect 528780 5842 528836 5852
rect 525196 4610 525252 4620
rect 529228 5796 529284 5806
rect 525420 4340 525476 4350
rect 525420 480 525476 4284
rect 527324 4228 527380 4238
rect 527324 480 527380 4172
rect 529228 480 529284 5740
rect 530572 4564 530628 8120
rect 530572 4498 530628 4508
rect 531132 6580 531188 6590
rect 531132 480 531188 6524
rect 532364 6580 532420 8120
rect 532364 6514 532420 6524
rect 533036 6692 533092 6702
rect 533036 480 533092 6636
rect 534156 4900 534212 8120
rect 534156 4834 534212 4844
rect 534940 6468 534996 6478
rect 534940 480 534996 6412
rect 535948 4452 536004 8120
rect 535948 4386 536004 4396
rect 536844 6356 536900 6366
rect 536844 480 536900 6300
rect 537740 4228 537796 8120
rect 539532 6468 539588 8120
rect 539532 6402 539588 6412
rect 537740 4162 537796 4172
rect 538748 6244 538804 6254
rect 538748 480 538804 6188
rect 540652 6132 540708 6142
rect 540652 480 540708 6076
rect 541324 4340 541380 8120
rect 543116 6356 543172 8120
rect 543116 6290 543172 6300
rect 544908 6244 544964 8120
rect 544908 6178 544964 6188
rect 546700 6132 546756 8120
rect 546700 6066 546756 6076
rect 544460 6020 544516 6030
rect 541324 4274 541380 4284
rect 542668 4676 542724 4686
rect 542668 480 542724 4620
rect 544460 480 544516 5964
rect 548492 6020 548548 8120
rect 548492 5954 548548 5964
rect 550172 6580 550228 6590
rect 546364 5908 546420 5918
rect 546364 480 546420 5852
rect 548268 4564 548324 4574
rect 548268 480 548324 4508
rect 550172 480 550228 6524
rect 550284 5908 550340 8120
rect 550284 5842 550340 5852
rect 552076 4676 552132 8120
rect 552076 4610 552132 4620
rect 552188 4900 552244 4910
rect 552188 480 552244 4844
rect 553868 4788 553924 8120
rect 553868 4722 553924 4732
rect 555660 4564 555716 8120
rect 557452 6580 557508 8120
rect 557452 6514 557508 6524
rect 555660 4498 555716 4508
rect 557788 6468 557844 6478
rect 553980 4452 554036 4462
rect 553980 480 554036 4396
rect 555884 4228 555940 4238
rect 555884 480 555940 4172
rect 557788 480 557844 6412
rect 559244 4228 559300 8120
rect 561036 6468 561092 8120
rect 561036 6402 561092 6412
rect 561596 6356 561652 6366
rect 559244 4162 559300 4172
rect 559692 4340 559748 4350
rect 559692 480 559748 4284
rect 561596 480 561652 6300
rect 562828 4452 562884 8120
rect 562828 4386 562884 4396
rect 563500 6244 563556 6254
rect 563500 480 563556 6188
rect 564620 4340 564676 8120
rect 564620 4274 564676 4284
rect 565404 6132 565460 6142
rect 565404 480 565460 6076
rect 567308 6020 567364 6030
rect 567308 480 567364 5964
rect 569212 5908 569268 5918
rect 569212 480 569268 5852
rect 573020 4788 573076 4798
rect 571228 4676 571284 4686
rect 571228 480 571284 4620
rect 573020 480 573076 4732
rect 574924 4564 574980 4574
rect 574924 480 574980 4508
rect 582540 4452 582596 4462
rect 578732 4228 578788 4238
rect 576828 3444 576884 3454
rect 576828 480 576884 3388
rect 578732 480 578788 4172
rect 580636 3444 580692 3454
rect 580636 480 580692 3388
rect 582540 480 582596 4396
rect 584444 4340 584500 4350
rect 584444 480 584500 4284
rect 270172 476 270536 480
rect 270172 420 270228 476
rect 269612 364 270228 420
rect 270284 392 270536 476
rect 272188 392 272440 480
rect 274092 392 274344 480
rect 275996 392 276248 480
rect 277900 392 278152 480
rect 279804 392 280056 480
rect 281708 392 281960 480
rect 283612 392 283864 480
rect 270312 -960 270536 392
rect 272216 -960 272440 392
rect 274120 -960 274344 392
rect 276024 -960 276248 392
rect 277928 -960 278152 392
rect 279832 -960 280056 392
rect 281736 -960 281960 392
rect 283640 -960 283864 392
rect 285544 -960 285768 480
rect 287420 392 287672 480
rect 289324 392 289576 480
rect 291228 392 291480 480
rect 293132 392 293384 480
rect 295036 392 295288 480
rect 296940 392 297192 480
rect 298844 392 299096 480
rect 300748 392 301000 480
rect 302652 392 302904 480
rect 304556 392 304808 480
rect 306460 392 306712 480
rect 308364 392 308616 480
rect 310268 392 310520 480
rect 312172 392 312424 480
rect 287448 -960 287672 392
rect 289352 -960 289576 392
rect 291256 -960 291480 392
rect 293160 -960 293384 392
rect 295064 -960 295288 392
rect 296968 -960 297192 392
rect 298872 -960 299096 392
rect 300776 -960 301000 392
rect 302680 -960 302904 392
rect 304584 -960 304808 392
rect 306488 -960 306712 392
rect 308392 -960 308616 392
rect 310296 -960 310520 392
rect 312200 -960 312424 392
rect 314104 -960 314328 480
rect 315980 392 316232 480
rect 317884 392 318136 480
rect 319788 392 320040 480
rect 321692 392 321944 480
rect 323596 392 323848 480
rect 325500 392 325752 480
rect 327404 392 327656 480
rect 329308 392 329560 480
rect 331212 392 331464 480
rect 333116 392 333368 480
rect 335020 392 335272 480
rect 336924 392 337176 480
rect 338828 392 339080 480
rect 340732 392 340984 480
rect 316008 -960 316232 392
rect 317912 -960 318136 392
rect 319816 -960 320040 392
rect 321720 -960 321944 392
rect 323624 -960 323848 392
rect 325528 -960 325752 392
rect 327432 -960 327656 392
rect 329336 -960 329560 392
rect 331240 -960 331464 392
rect 333144 -960 333368 392
rect 335048 -960 335272 392
rect 336952 -960 337176 392
rect 338856 -960 339080 392
rect 340760 -960 340984 392
rect 342664 -960 342888 480
rect 344540 392 344792 480
rect 346444 392 346696 480
rect 348348 392 348600 480
rect 350252 392 350504 480
rect 352156 392 352408 480
rect 354060 392 354312 480
rect 355964 392 356216 480
rect 357868 392 358120 480
rect 359772 392 360024 480
rect 361676 392 361928 480
rect 363580 392 363832 480
rect 365484 392 365736 480
rect 367388 392 367640 480
rect 369292 392 369544 480
rect 344568 -960 344792 392
rect 346472 -960 346696 392
rect 348376 -960 348600 392
rect 350280 -960 350504 392
rect 352184 -960 352408 392
rect 354088 -960 354312 392
rect 355992 -960 356216 392
rect 357896 -960 358120 392
rect 359800 -960 360024 392
rect 361704 -960 361928 392
rect 363608 -960 363832 392
rect 365512 -960 365736 392
rect 367416 -960 367640 392
rect 369320 -960 369544 392
rect 371224 -960 371448 480
rect 373100 392 373352 480
rect 375004 392 375256 480
rect 376908 392 377160 480
rect 378812 392 379064 480
rect 380716 392 380968 480
rect 382620 392 382872 480
rect 384524 392 384776 480
rect 386428 392 386680 480
rect 388332 392 388584 480
rect 390236 392 390488 480
rect 392140 392 392392 480
rect 394044 392 394296 480
rect 395948 392 396200 480
rect 397852 392 398104 480
rect 373128 -960 373352 392
rect 375032 -960 375256 392
rect 376936 -960 377160 392
rect 378840 -960 379064 392
rect 380744 -960 380968 392
rect 382648 -960 382872 392
rect 384552 -960 384776 392
rect 386456 -960 386680 392
rect 388360 -960 388584 392
rect 390264 -960 390488 392
rect 392168 -960 392392 392
rect 394072 -960 394296 392
rect 395976 -960 396200 392
rect 397880 -960 398104 392
rect 399784 -960 400008 480
rect 401660 392 401912 480
rect 403564 392 403816 480
rect 405468 392 405720 480
rect 407372 392 407624 480
rect 409276 392 409528 480
rect 411180 392 411432 480
rect 413084 392 413336 480
rect 414988 392 415240 480
rect 416892 392 417144 480
rect 418796 392 419048 480
rect 420700 392 420952 480
rect 422604 392 422856 480
rect 424508 392 424760 480
rect 426412 392 426664 480
rect 401688 -960 401912 392
rect 403592 -960 403816 392
rect 405496 -960 405720 392
rect 407400 -960 407624 392
rect 409304 -960 409528 392
rect 411208 -960 411432 392
rect 413112 -960 413336 392
rect 415016 -960 415240 392
rect 416920 -960 417144 392
rect 418824 -960 419048 392
rect 420728 -960 420952 392
rect 422632 -960 422856 392
rect 424536 -960 424760 392
rect 426440 -960 426664 392
rect 428344 -960 428568 480
rect 430248 -960 430472 480
rect 432124 392 432376 480
rect 434028 392 434280 480
rect 435932 392 436184 480
rect 437836 392 438088 480
rect 439740 392 439992 480
rect 441644 392 441896 480
rect 443548 392 443800 480
rect 445452 392 445704 480
rect 447356 392 447608 480
rect 449260 392 449512 480
rect 451164 392 451416 480
rect 453068 392 453320 480
rect 454972 392 455224 480
rect 432152 -960 432376 392
rect 434056 -960 434280 392
rect 435960 -960 436184 392
rect 437864 -960 438088 392
rect 439768 -960 439992 392
rect 441672 -960 441896 392
rect 443576 -960 443800 392
rect 445480 -960 445704 392
rect 447384 -960 447608 392
rect 449288 -960 449512 392
rect 451192 -960 451416 392
rect 453096 -960 453320 392
rect 455000 -960 455224 392
rect 456904 -960 457128 480
rect 458780 392 459032 480
rect 460684 392 460936 480
rect 462588 392 462840 480
rect 464492 392 464744 480
rect 466396 392 466648 480
rect 468300 392 468552 480
rect 470204 392 470456 480
rect 472108 392 472360 480
rect 474012 392 474264 480
rect 475916 392 476168 480
rect 477820 392 478072 480
rect 479724 392 479976 480
rect 481628 392 481880 480
rect 483532 392 483784 480
rect 458808 -960 459032 392
rect 460712 -960 460936 392
rect 462616 -960 462840 392
rect 464520 -960 464744 392
rect 466424 -960 466648 392
rect 468328 -960 468552 392
rect 470232 -960 470456 392
rect 472136 -960 472360 392
rect 474040 -960 474264 392
rect 475944 -960 476168 392
rect 477848 -960 478072 392
rect 479752 -960 479976 392
rect 481656 -960 481880 392
rect 483560 -960 483784 392
rect 485464 -960 485688 480
rect 487340 392 487592 480
rect 489244 392 489496 480
rect 491148 392 491400 480
rect 493052 392 493304 480
rect 494956 392 495208 480
rect 496860 392 497112 480
rect 498764 392 499016 480
rect 500668 392 500920 480
rect 502572 392 502824 480
rect 504476 392 504728 480
rect 506380 392 506632 480
rect 508284 392 508536 480
rect 510188 392 510440 480
rect 512092 392 512344 480
rect 487368 -960 487592 392
rect 489272 -960 489496 392
rect 491176 -960 491400 392
rect 493080 -960 493304 392
rect 494984 -960 495208 392
rect 496888 -960 497112 392
rect 498792 -960 499016 392
rect 500696 -960 500920 392
rect 502600 -960 502824 392
rect 504504 -960 504728 392
rect 506408 -960 506632 392
rect 508312 -960 508536 392
rect 510216 -960 510440 392
rect 512120 -960 512344 392
rect 514024 -960 514248 480
rect 515900 392 516152 480
rect 517804 392 518056 480
rect 519708 392 519960 480
rect 521612 392 521864 480
rect 523516 392 523768 480
rect 525420 392 525672 480
rect 527324 392 527576 480
rect 529228 392 529480 480
rect 531132 392 531384 480
rect 533036 392 533288 480
rect 534940 392 535192 480
rect 536844 392 537096 480
rect 538748 392 539000 480
rect 540652 392 540904 480
rect 515928 -960 516152 392
rect 517832 -960 518056 392
rect 519736 -960 519960 392
rect 521640 -960 521864 392
rect 523544 -960 523768 392
rect 525448 -960 525672 392
rect 527352 -960 527576 392
rect 529256 -960 529480 392
rect 531160 -960 531384 392
rect 533064 -960 533288 392
rect 534968 -960 535192 392
rect 536872 -960 537096 392
rect 538776 -960 539000 392
rect 540680 -960 540904 392
rect 542584 -960 542808 480
rect 544460 392 544712 480
rect 546364 392 546616 480
rect 548268 392 548520 480
rect 550172 392 550424 480
rect 544488 -960 544712 392
rect 546392 -960 546616 392
rect 548296 -960 548520 392
rect 550200 -960 550424 392
rect 552104 -960 552328 480
rect 553980 392 554232 480
rect 555884 392 556136 480
rect 557788 392 558040 480
rect 559692 392 559944 480
rect 561596 392 561848 480
rect 563500 392 563752 480
rect 565404 392 565656 480
rect 567308 392 567560 480
rect 569212 392 569464 480
rect 554008 -960 554232 392
rect 555912 -960 556136 392
rect 557816 -960 558040 392
rect 559720 -960 559944 392
rect 561624 -960 561848 392
rect 563528 -960 563752 392
rect 565432 -960 565656 392
rect 567336 -960 567560 392
rect 569240 -960 569464 392
rect 571144 -960 571368 480
rect 573020 392 573272 480
rect 574924 392 575176 480
rect 576828 392 577080 480
rect 578732 392 578984 480
rect 580636 392 580888 480
rect 582540 392 582792 480
rect 584444 392 584696 480
rect 573048 -960 573272 392
rect 574952 -960 575176 392
rect 576856 -960 577080 392
rect 578760 -960 578984 392
rect 580664 -960 580888 392
rect 582568 -960 582792 392
rect 584472 -960 584696 392
<< via2 >>
rect 11228 588812 11284 588868
rect 16492 588812 16548 588868
rect 48300 591276 48356 591332
rect 55132 591276 55188 591332
rect 77420 591276 77476 591332
rect 80108 591276 80164 591332
rect 96012 591276 96068 591332
rect 99260 591276 99316 591332
rect 111916 588812 111972 588868
rect 121324 588812 121380 588868
rect 159628 590492 159684 590548
rect 165452 590492 165508 590548
rect 175532 588812 175588 588868
rect 187516 588812 187572 588868
rect 207340 591276 207396 591332
rect 209580 591276 209636 591332
rect 223244 590492 223300 590548
rect 231644 590492 231700 590548
rect 239148 588812 239204 588868
rect 253708 588812 253764 588868
rect 270956 591276 271012 591332
rect 275772 591276 275828 591332
rect 286860 588812 286916 588868
rect 297836 588812 297892 588868
rect 302764 588812 302820 588868
rect 319900 588812 319956 588868
rect 334572 590492 334628 590548
rect 341964 590492 342020 590548
rect 350476 590492 350532 590548
rect 364028 590492 364084 590548
rect 366380 588812 366436 588868
rect 386092 588812 386148 588868
rect 398188 588812 398244 588868
rect 429996 590492 430052 590548
rect 408268 588812 408324 588868
rect 414092 588812 414148 588868
rect 452284 590492 452340 590548
rect 461804 590492 461860 590548
rect 430220 588812 430276 588868
rect 474348 590492 474404 590548
rect 493612 590492 493668 590548
rect 477708 588812 477764 588868
rect 518476 590492 518532 590548
rect 496412 588812 496468 588868
rect 525420 588812 525476 588868
rect 540540 588812 540596 588868
rect 541324 590604 541380 590660
rect 562604 590604 562660 590660
rect 557228 590492 557284 590548
rect 584668 590492 584724 590548
rect 11564 5852 11620 5908
rect 25228 5852 25284 5908
rect 26796 4956 26852 5012
rect 24892 4844 24948 4900
rect 22988 4732 23044 4788
rect 21084 4620 21140 4676
rect 19180 4508 19236 4564
rect 17276 4396 17332 4452
rect 15372 4284 15428 4340
rect 13356 4172 13412 4228
rect 39564 4956 39620 5012
rect 37772 4844 37828 4900
rect 35980 4732 36036 4788
rect 40124 4732 40180 4788
rect 34188 4620 34244 4676
rect 38220 4620 38276 4676
rect 32396 4508 32452 4564
rect 36316 4508 36372 4564
rect 30604 4396 30660 4452
rect 34412 4396 34468 4452
rect 28812 4284 28868 4340
rect 32508 4284 32564 4340
rect 27020 4172 27076 4228
rect 30604 4172 30660 4228
rect 28700 4060 28756 4116
rect 41356 4060 41412 4116
rect 41916 4844 41972 4900
rect 53900 4844 53956 4900
rect 55356 4844 55412 4900
rect 52108 4732 52164 4788
rect 53452 4732 53508 4788
rect 50316 4620 50372 4676
rect 51548 4620 51604 4676
rect 48524 4508 48580 4564
rect 49644 4508 49700 4564
rect 46732 4396 46788 4452
rect 47740 4396 47796 4452
rect 44940 4284 44996 4340
rect 45836 4284 45892 4340
rect 43148 4172 43204 4228
rect 43932 4172 43988 4228
rect 64652 4732 64708 4788
rect 64876 4956 64932 5012
rect 62860 4620 62916 4676
rect 61068 4508 61124 4564
rect 62972 4508 63028 4564
rect 59276 4396 59332 4452
rect 61180 4396 61236 4452
rect 57484 4284 57540 4340
rect 55692 4172 55748 4228
rect 57260 4172 57316 4228
rect 59164 4060 59220 4116
rect 66444 4844 66500 4900
rect 66780 4620 66836 4676
rect 68236 4172 68292 4228
rect 68684 4172 68740 4228
rect 75404 4956 75460 5012
rect 76300 4732 76356 4788
rect 73612 4508 73668 4564
rect 74396 4508 74452 4564
rect 71820 4396 71876 4452
rect 72492 4396 72548 4452
rect 70028 4060 70084 4116
rect 70476 4284 70532 4340
rect 77196 4620 77252 4676
rect 78204 4620 78260 4676
rect 86156 4732 86212 4788
rect 87724 4732 87780 4788
rect 84364 4508 84420 4564
rect 85820 4508 85876 4564
rect 82572 4396 82628 4452
rect 80780 4284 80836 4340
rect 82012 4284 82068 4340
rect 78988 4172 79044 4228
rect 80108 4172 80164 4228
rect 83916 4060 83972 4116
rect 87948 4620 88004 4676
rect 89628 4620 89684 4676
rect 90860 4284 90916 4340
rect 89740 4172 89796 4228
rect 91532 4172 91588 4228
rect 96908 4732 96964 4788
rect 98700 4620 98756 4676
rect 95116 4508 95172 4564
rect 99036 4508 99092 4564
rect 97244 4396 97300 4452
rect 93324 4060 93380 4116
rect 93436 4284 93492 4340
rect 95340 4060 95396 4116
rect 102284 4284 102340 4340
rect 102956 4284 103012 4340
rect 100492 4172 100548 4228
rect 101052 4172 101108 4228
rect 104076 4060 104132 4116
rect 104860 4620 104916 4676
rect 107660 4508 107716 4564
rect 105868 4396 105924 4452
rect 113036 4620 113092 4676
rect 114380 4620 114436 4676
rect 111244 4284 111300 4340
rect 112476 4284 112532 4340
rect 109452 4172 109508 4228
rect 110572 4172 110628 4228
rect 108668 4060 108724 4116
rect 106764 3948 106820 4004
rect 114828 3948 114884 4004
rect 116284 4396 116340 4452
rect 121996 4620 122052 4676
rect 123788 4396 123844 4452
rect 123900 4620 123956 4676
rect 120204 4284 120260 4340
rect 118412 4172 118468 4228
rect 116620 4060 116676 4116
rect 121996 4060 122052 4116
rect 120092 3948 120148 4004
rect 118188 3836 118244 3892
rect 125580 3836 125636 3892
rect 125804 4732 125860 4788
rect 127372 3948 127428 4004
rect 127596 4396 127652 4452
rect 132748 4732 132804 4788
rect 130956 4620 131012 4676
rect 134540 4396 134596 4452
rect 135324 4396 135380 4452
rect 129164 4060 129220 4116
rect 129612 4172 129668 4228
rect 133420 4060 133476 4116
rect 131516 3948 131572 4004
rect 136332 4172 136388 4228
rect 137228 4172 137284 4228
rect 138124 3948 138180 4004
rect 139132 4284 139188 4340
rect 139916 4060 139972 4116
rect 141036 4508 141092 4564
rect 141708 4396 141764 4452
rect 145292 4284 145348 4340
rect 146748 4620 146804 4676
rect 143500 4172 143556 4228
rect 144844 4060 144900 4116
rect 142940 3948 142996 4004
rect 147084 4508 147140 4564
rect 148652 4508 148708 4564
rect 148876 3948 148932 4004
rect 150556 4396 150612 4452
rect 152460 4620 152516 4676
rect 154252 4508 154308 4564
rect 156044 4396 156100 4452
rect 150668 4060 150724 4116
rect 152460 4172 152516 4228
rect 157836 4172 157892 4228
rect 158172 4060 158228 4116
rect 156156 3948 156212 4004
rect 154364 3836 154420 3892
rect 159628 3836 159684 3892
rect 160076 4172 160132 4228
rect 161420 3948 161476 4004
rect 161980 4284 162036 4340
rect 163212 4060 163268 4116
rect 163884 4396 163940 4452
rect 168588 4396 168644 4452
rect 166796 4284 166852 4340
rect 165004 4172 165060 4228
rect 165788 4172 165844 4228
rect 170380 4172 170436 4228
rect 171500 5068 171556 5124
rect 169596 4060 169652 4116
rect 167692 3948 167748 4004
rect 172172 3948 172228 4004
rect 173404 5964 173460 6020
rect 173964 4060 174020 4116
rect 175308 6076 175364 6132
rect 179340 6076 179396 6132
rect 177548 5964 177604 6020
rect 175756 5068 175812 5124
rect 177212 5292 177268 5348
rect 181132 5292 181188 5348
rect 179116 5180 179172 5236
rect 182924 5180 182980 5236
rect 181020 5068 181076 5124
rect 184716 5068 184772 5124
rect 184716 4284 184772 4340
rect 182924 4060 182980 4116
rect 186508 4060 186564 4116
rect 186732 5852 186788 5908
rect 190092 5852 190148 5908
rect 190540 5180 190596 5236
rect 188300 4284 188356 4340
rect 188636 5068 188692 5124
rect 193676 5180 193732 5236
rect 194348 5180 194404 5236
rect 191884 5068 191940 5124
rect 192444 5068 192500 5124
rect 197260 5180 197316 5236
rect 198156 5852 198212 5908
rect 195468 5068 195524 5124
rect 196252 5068 196308 5124
rect 200844 5852 200900 5908
rect 199052 5068 199108 5124
rect 200060 5180 200116 5236
rect 202636 5180 202692 5236
rect 203868 5180 203924 5236
rect 201964 5068 202020 5124
rect 206220 5180 206276 5236
rect 207676 5180 207732 5236
rect 204428 5068 204484 5124
rect 205772 5068 205828 5124
rect 209804 5180 209860 5236
rect 211484 5964 211540 6020
rect 208012 5068 208068 5124
rect 209580 5068 209636 5124
rect 213388 5964 213444 6020
rect 211596 5068 211652 5124
rect 213276 5180 213332 5236
rect 215180 5180 215236 5236
rect 215292 5068 215348 5124
rect 216972 5068 217028 5124
rect 217196 5068 217252 5124
rect 218764 5068 218820 5124
rect 222908 5852 222964 5908
rect 224140 5852 224196 5908
rect 258188 5852 258244 5908
rect 258860 5852 258916 5908
rect 265356 5068 265412 5124
rect 266476 5068 266532 5124
rect 270732 5068 270788 5124
rect 272188 5068 272244 5124
rect 272524 5068 272580 5124
rect 274092 5068 274148 5124
rect 277900 5404 277956 5460
rect 276108 5180 276164 5236
rect 277900 5180 277956 5236
rect 274316 5068 274372 5124
rect 275996 5068 276052 5124
rect 281484 5852 281540 5908
rect 279692 5068 279748 5124
rect 279804 5404 279860 5460
rect 281708 5068 281764 5124
rect 283276 4060 283332 4116
rect 283612 5852 283668 5908
rect 285068 3948 285124 4004
rect 285628 4060 285684 4116
rect 286860 4060 286916 4116
rect 287420 3948 287476 4004
rect 288652 3948 288708 4004
rect 289324 4060 289380 4116
rect 295820 5180 295876 5236
rect 294028 5068 294084 5124
rect 296940 5068 296996 5124
rect 292236 4172 292292 4228
rect 295036 4172 295092 4228
rect 290444 4060 290500 4116
rect 293132 4060 293188 4116
rect 291228 3948 291284 4004
rect 297612 4060 297668 4116
rect 298844 5180 298900 5236
rect 299404 3948 299460 4004
rect 300748 4060 300804 4116
rect 304780 4396 304836 4452
rect 302988 4172 303044 4228
rect 306460 4172 306516 4228
rect 301196 4060 301252 4116
rect 304556 4060 304612 4116
rect 302652 3948 302708 4004
rect 315532 6076 315588 6132
rect 317324 5964 317380 6020
rect 313740 5852 313796 5908
rect 317884 5852 317940 5908
rect 311948 5180 312004 5236
rect 315980 5180 316036 5236
rect 310156 5068 310212 5124
rect 314188 5068 314244 5124
rect 308364 4620 308420 4676
rect 312172 4620 312228 4676
rect 306572 4060 306628 4116
rect 308364 4396 308420 4452
rect 310268 4060 310324 4116
rect 319116 5068 319172 5124
rect 319788 6076 319844 6132
rect 320908 4060 320964 4116
rect 321692 5964 321748 6020
rect 324492 5964 324548 6020
rect 328076 6076 328132 6132
rect 326284 5852 326340 5908
rect 329308 5964 329364 6020
rect 322700 3948 322756 4004
rect 323596 5068 323652 5124
rect 325500 4060 325556 4116
rect 327404 3948 327460 4004
rect 329868 5068 329924 5124
rect 331212 5852 331268 5908
rect 331660 5180 331716 5236
rect 333116 6076 333172 6132
rect 333452 5292 333508 5348
rect 335020 5068 335076 5124
rect 337036 6076 337092 6132
rect 338828 5964 338884 6020
rect 340620 5852 340676 5908
rect 338828 5292 338884 5348
rect 335244 5068 335300 5124
rect 336924 5180 336980 5236
rect 340732 5068 340788 5124
rect 342412 5068 342468 5124
rect 342748 6076 342804 6132
rect 344204 5180 344260 5236
rect 344540 5964 344596 6020
rect 345996 5292 346052 5348
rect 346444 5852 346500 5908
rect 349580 6188 349636 6244
rect 351372 6076 351428 6132
rect 347788 5852 347844 5908
rect 352156 5292 352212 5348
rect 350252 5180 350308 5236
rect 348348 5068 348404 5124
rect 353164 5068 353220 5124
rect 354060 5852 354116 5908
rect 354956 5180 355012 5236
rect 355964 6188 356020 6244
rect 356748 5292 356804 5348
rect 357868 6076 357924 6132
rect 358540 6076 358596 6132
rect 360332 5964 360388 6020
rect 362124 5852 362180 5908
rect 363580 5292 363636 5348
rect 361676 5180 361732 5236
rect 359772 5068 359828 5124
rect 363916 4396 363972 4452
rect 365484 6076 365540 6132
rect 365708 4060 365764 4116
rect 367388 5964 367444 6020
rect 367500 3948 367556 4004
rect 369292 5852 369348 5908
rect 369516 4284 369572 4340
rect 371084 4172 371140 4228
rect 371308 4396 371364 4452
rect 374668 5964 374724 6020
rect 376460 5068 376516 5124
rect 372876 4396 372932 4452
rect 376908 4284 376964 4340
rect 373100 4060 373156 4116
rect 375004 3948 375060 4004
rect 378252 4060 378308 4116
rect 378812 4172 378868 4228
rect 381836 4620 381892 4676
rect 382620 5964 382676 6020
rect 380044 4172 380100 4228
rect 380716 4396 380772 4452
rect 383628 4508 383684 4564
rect 384524 5068 384580 5124
rect 385420 4396 385476 4452
rect 387212 4284 387268 4340
rect 388332 4172 388388 4228
rect 386428 4060 386484 4116
rect 392588 6412 392644 6468
rect 390796 6300 390852 6356
rect 396172 6188 396228 6244
rect 397964 6076 398020 6132
rect 399756 5964 399812 6020
rect 399868 6300 399924 6356
rect 394380 5852 394436 5908
rect 389004 4060 389060 4116
rect 390236 4620 390292 4676
rect 392140 4508 392196 4564
rect 394044 4396 394100 4452
rect 395948 4284 396004 4340
rect 397852 4060 397908 4116
rect 401548 4060 401604 4116
rect 401660 6412 401716 6468
rect 403340 4172 403396 4228
rect 403564 5852 403620 5908
rect 408716 6412 408772 6468
rect 406924 6300 406980 6356
rect 405132 5852 405188 5908
rect 405468 6188 405524 6244
rect 410508 6188 410564 6244
rect 407372 6076 407428 6132
rect 409276 5964 409332 6020
rect 414092 5964 414148 6020
rect 412300 5068 412356 5124
rect 414988 5852 415044 5908
rect 413084 4172 413140 4228
rect 411180 4060 411236 4116
rect 415884 5852 415940 5908
rect 416892 6300 416948 6356
rect 419468 6636 419524 6692
rect 417676 6300 417732 6356
rect 418796 6412 418852 6468
rect 423052 6524 423108 6580
rect 421260 6412 421316 6468
rect 420700 6188 420756 6244
rect 424844 6188 424900 6244
rect 426636 6076 426692 6132
rect 428428 6300 428484 6356
rect 424508 5964 424564 6020
rect 422604 5068 422660 5124
rect 426412 5852 426468 5908
rect 429100 5964 429156 6020
rect 430220 5852 430276 5908
rect 430332 6636 430388 6692
rect 432012 6300 432068 6356
rect 432124 6412 432180 6468
rect 433804 6412 433860 6468
rect 434028 6524 434084 6580
rect 435596 6524 435652 6580
rect 435932 6188 435988 6244
rect 437388 6188 437444 6244
rect 437836 6076 437892 6132
rect 439180 6076 439236 6132
rect 439740 5964 439796 6020
rect 440972 5964 441028 6020
rect 441644 5852 441700 5908
rect 442764 5852 442820 5908
rect 443548 6300 443604 6356
rect 444556 6300 444612 6356
rect 445452 6412 445508 6468
rect 446348 6412 446404 6468
rect 447356 6524 447412 6580
rect 448140 5740 448196 5796
rect 449260 6188 449316 6244
rect 449932 6188 449988 6244
rect 451164 6076 451220 6132
rect 451724 6076 451780 6132
rect 453068 5964 453124 6020
rect 453516 5964 453572 6020
rect 454972 5852 455028 5908
rect 457100 6636 457156 6692
rect 458892 6524 458948 6580
rect 458780 6412 458836 6468
rect 455308 5852 455364 5908
rect 456988 6300 457044 6356
rect 460684 6412 460740 6468
rect 462476 6300 462532 6356
rect 462588 6188 462644 6244
rect 460684 5740 460740 5796
rect 464268 6188 464324 6244
rect 464492 6076 464548 6132
rect 466060 6076 466116 6132
rect 466396 5964 466452 6020
rect 467852 5964 467908 6020
rect 468300 5852 468356 5908
rect 469644 5852 469700 5908
rect 470204 6636 470260 6692
rect 471436 4620 471492 4676
rect 472108 6524 472164 6580
rect 473228 4732 473284 4788
rect 474012 6412 474068 6468
rect 475020 4508 475076 4564
rect 475916 6300 475972 6356
rect 476812 4284 476868 4340
rect 477820 6188 477876 6244
rect 478604 4172 478660 4228
rect 479724 6076 479780 6132
rect 480396 4396 480452 4452
rect 481628 5964 481684 6020
rect 482188 5964 482244 6020
rect 483532 5852 483588 5908
rect 483980 5852 484036 5908
rect 485772 4844 485828 4900
rect 487340 4732 487396 4788
rect 485548 4620 485604 4676
rect 487564 4732 487620 4788
rect 489356 4620 489412 4676
rect 489244 4508 489300 4564
rect 491148 4508 491204 4564
rect 491148 4284 491204 4340
rect 492940 4284 492996 4340
rect 493052 4172 493108 4228
rect 494732 4172 494788 4228
rect 494956 4396 495012 4452
rect 500108 6412 500164 6468
rect 498316 6300 498372 6356
rect 501900 6188 501956 6244
rect 503692 6076 503748 6132
rect 496524 4396 496580 4452
rect 496860 5964 496916 6020
rect 505484 5964 505540 6020
rect 498764 5852 498820 5908
rect 507276 5852 507332 5908
rect 500668 4844 500724 4900
rect 502572 4732 502628 4788
rect 504476 4620 504532 4676
rect 506380 4508 506436 4564
rect 508284 4284 508340 4340
rect 509068 4284 509124 4340
rect 510188 4172 510244 4228
rect 516236 6636 516292 6692
rect 514444 6524 514500 6580
rect 515900 6412 515956 6468
rect 512652 5740 512708 5796
rect 514108 6300 514164 6356
rect 510860 4172 510916 4228
rect 512092 4396 512148 4452
rect 518028 6412 518084 6468
rect 519820 6300 519876 6356
rect 517804 6188 517860 6244
rect 521612 6188 521668 6244
rect 519708 6076 519764 6132
rect 523404 6076 523460 6132
rect 521612 5964 521668 6020
rect 523516 5852 523572 5908
rect 526988 5964 527044 6020
rect 528780 5852 528836 5908
rect 525196 4620 525252 4676
rect 529228 5740 529284 5796
rect 525420 4284 525476 4340
rect 527324 4172 527380 4228
rect 530572 4508 530628 4564
rect 531132 6524 531188 6580
rect 532364 6524 532420 6580
rect 533036 6636 533092 6692
rect 534156 4844 534212 4900
rect 534940 6412 534996 6468
rect 535948 4396 536004 4452
rect 536844 6300 536900 6356
rect 539532 6412 539588 6468
rect 537740 4172 537796 4228
rect 538748 6188 538804 6244
rect 540652 6076 540708 6132
rect 543116 6300 543172 6356
rect 544908 6188 544964 6244
rect 546700 6076 546756 6132
rect 544460 5964 544516 6020
rect 541324 4284 541380 4340
rect 542668 4620 542724 4676
rect 548492 5964 548548 6020
rect 550172 6524 550228 6580
rect 546364 5852 546420 5908
rect 548268 4508 548324 4564
rect 550284 5852 550340 5908
rect 552076 4620 552132 4676
rect 552188 4844 552244 4900
rect 553868 4732 553924 4788
rect 557452 6524 557508 6580
rect 555660 4508 555716 4564
rect 557788 6412 557844 6468
rect 553980 4396 554036 4452
rect 555884 4172 555940 4228
rect 561036 6412 561092 6468
rect 561596 6300 561652 6356
rect 559244 4172 559300 4228
rect 559692 4284 559748 4340
rect 562828 4396 562884 4452
rect 563500 6188 563556 6244
rect 564620 4284 564676 4340
rect 565404 6076 565460 6132
rect 567308 5964 567364 6020
rect 569212 5852 569268 5908
rect 573020 4732 573076 4788
rect 571228 4620 571284 4676
rect 574924 4508 574980 4564
rect 582540 4396 582596 4452
rect 578732 4172 578788 4228
rect 576828 3388 576884 3444
rect 580636 3388 580692 3444
rect 584444 4284 584500 4340
<< metal3 >>
rect 48290 591276 48300 591332
rect 48356 591276 55132 591332
rect 55188 591276 55198 591332
rect 77410 591276 77420 591332
rect 77476 591276 80108 591332
rect 80164 591276 80174 591332
rect 96002 591276 96012 591332
rect 96068 591276 99260 591332
rect 99316 591276 99326 591332
rect 207330 591276 207340 591332
rect 207396 591276 209580 591332
rect 209636 591276 209646 591332
rect 270946 591276 270956 591332
rect 271012 591276 275772 591332
rect 275828 591276 275838 591332
rect 541314 590604 541324 590660
rect 541380 590604 562604 590660
rect 562660 590604 562670 590660
rect 159618 590492 159628 590548
rect 159684 590492 165452 590548
rect 165508 590492 165518 590548
rect 223234 590492 223244 590548
rect 223300 590492 231644 590548
rect 231700 590492 231710 590548
rect 334562 590492 334572 590548
rect 334628 590492 341964 590548
rect 342020 590492 342030 590548
rect 350466 590492 350476 590548
rect 350532 590492 364028 590548
rect 364084 590492 364094 590548
rect 429986 590492 429996 590548
rect 430052 590492 452284 590548
rect 452340 590492 452350 590548
rect 461794 590492 461804 590548
rect 461860 590492 474348 590548
rect 474404 590492 474414 590548
rect 493602 590492 493612 590548
rect 493668 590492 518476 590548
rect 518532 590492 518542 590548
rect 557218 590492 557228 590548
rect 557284 590492 584668 590548
rect 584724 590492 584734 590548
rect 11218 588812 11228 588868
rect 11284 588812 16492 588868
rect 16548 588812 16558 588868
rect 111906 588812 111916 588868
rect 111972 588812 121324 588868
rect 121380 588812 121390 588868
rect 175522 588812 175532 588868
rect 175588 588812 187516 588868
rect 187572 588812 187582 588868
rect 239138 588812 239148 588868
rect 239204 588812 253708 588868
rect 253764 588812 253774 588868
rect 286850 588812 286860 588868
rect 286916 588812 297836 588868
rect 297892 588812 297902 588868
rect 302754 588812 302764 588868
rect 302820 588812 319900 588868
rect 319956 588812 319966 588868
rect 366370 588812 366380 588868
rect 366436 588812 386092 588868
rect 386148 588812 386158 588868
rect 398178 588812 398188 588868
rect 398244 588812 408268 588868
rect 408324 588812 408334 588868
rect 414082 588812 414092 588868
rect 414148 588812 430220 588868
rect 430276 588812 430286 588868
rect 477698 588812 477708 588868
rect 477764 588812 496412 588868
rect 496468 588812 496478 588868
rect 525410 588812 525420 588868
rect 525476 588812 540540 588868
rect 540596 588812 540606 588868
rect 595560 588644 597000 588840
rect 590482 588588 590492 588644
rect 590548 588616 597000 588644
rect 590548 588588 595672 588616
rect -960 587188 480 587384
rect -960 587160 4172 587188
rect 392 587132 4172 587160
rect 4228 587132 4238 587188
rect 582008 576268 590492 576324
rect 590548 576268 590558 576324
rect 595560 575428 597000 575624
rect 591266 575372 591276 575428
rect 591332 575400 597000 575428
rect 591332 575372 595672 575400
rect -960 573076 480 573272
rect -960 573048 4284 573076
rect 392 573020 4284 573048
rect 4340 573020 4350 573076
rect 582008 565516 591276 565572
rect 591332 565516 591342 565572
rect 4162 565068 4172 565124
rect 4228 565068 8120 565124
rect 595560 562212 597000 562408
rect 586338 562156 586348 562212
rect 586404 562184 597000 562212
rect 586404 562156 595672 562184
rect -960 558964 480 559160
rect -960 558936 6188 558964
rect 392 558908 6188 558936
rect 6244 558908 6254 558964
rect 582008 554764 586348 554820
rect 586404 554764 586414 554820
rect 4274 554540 4284 554596
rect 4340 554540 8120 554596
rect 595560 548996 597000 549192
rect 590482 548940 590492 548996
rect 590548 548968 597000 548996
rect 590548 548940 595672 548968
rect -960 544852 480 545048
rect -960 544824 4172 544852
rect 392 544796 4172 544824
rect 4228 544796 4238 544852
rect 6178 544012 6188 544068
rect 6244 544012 8120 544068
rect 595560 535780 597000 535976
rect 588578 535724 588588 535780
rect 588644 535752 597000 535780
rect 588644 535724 595672 535752
rect 582008 533260 590492 533316
rect 590548 533260 590558 533316
rect -960 530740 480 530936
rect -960 530712 4284 530740
rect 392 530684 4284 530712
rect 4340 530684 4350 530740
rect 4162 522956 4172 523012
rect 4228 522956 8120 523012
rect 595560 522564 597000 522760
rect 582008 522508 588588 522564
rect 588644 522508 588654 522564
rect 588802 522508 588812 522564
rect 588868 522536 597000 522564
rect 588868 522508 595672 522536
rect -960 516628 480 516824
rect -960 516600 6188 516628
rect 392 516572 6188 516600
rect 6244 516572 6254 516628
rect 4274 512428 4284 512484
rect 4340 512428 8120 512484
rect 582008 511756 588812 511812
rect 588868 511756 588878 511812
rect 595560 509348 597000 509544
rect 585442 509292 585452 509348
rect 585508 509320 597000 509348
rect 585508 509292 595672 509320
rect -960 502516 480 502712
rect -960 502488 4172 502516
rect 392 502460 4172 502488
rect 4228 502460 4238 502516
rect 6178 501900 6188 501956
rect 6244 501900 8120 501956
rect 595560 496132 597000 496328
rect 590482 496076 590492 496132
rect 590548 496104 597000 496132
rect 590548 496076 595672 496104
rect 582008 490252 585452 490308
rect 585508 490252 585518 490308
rect -960 488404 480 488600
rect -960 488376 4284 488404
rect 392 488348 4284 488376
rect 4340 488348 4350 488404
rect 595560 482916 597000 483112
rect 590594 482860 590604 482916
rect 590660 482888 597000 482916
rect 590660 482860 595672 482888
rect 4162 480844 4172 480900
rect 4228 480844 8120 480900
rect 582008 479500 590492 479556
rect 590548 479500 590558 479556
rect -960 474292 480 474488
rect -960 474264 6412 474292
rect 392 474236 6412 474264
rect 6468 474236 6478 474292
rect 4274 470316 4284 470372
rect 4340 470316 8120 470372
rect 595560 469700 597000 469896
rect 585442 469644 585452 469700
rect 585508 469672 597000 469700
rect 585508 469644 595672 469672
rect 582008 468748 590604 468804
rect 590660 468748 590670 468804
rect -960 460180 480 460376
rect -960 460152 6188 460180
rect 392 460124 6188 460152
rect 6244 460124 6254 460180
rect 6402 459788 6412 459844
rect 6468 459788 8120 459844
rect 595560 456484 597000 456680
rect 585554 456428 585564 456484
rect 585620 456456 597000 456484
rect 585620 456428 595672 456456
rect 582008 447244 585452 447300
rect 585508 447244 585518 447300
rect -960 446068 480 446264
rect -960 446040 4172 446068
rect 392 446012 4172 446040
rect 4228 446012 4238 446068
rect 595560 443268 597000 443464
rect 590482 443212 590492 443268
rect 590548 443240 597000 443268
rect 590548 443212 595672 443240
rect 6178 438732 6188 438788
rect 6244 438732 8120 438788
rect 582008 436492 585564 436548
rect 585620 436492 585630 436548
rect -960 431956 480 432152
rect -960 431928 6412 431956
rect 392 431900 6412 431928
rect 6468 431900 6478 431956
rect 595560 430164 597000 430248
rect 585442 430108 585452 430164
rect 585508 430108 597000 430164
rect 595560 430024 597000 430108
rect 4162 428204 4172 428260
rect 4228 428204 8120 428260
rect 582008 425740 590492 425796
rect 590548 425740 590558 425796
rect -960 417844 480 418040
rect -960 417816 6188 417844
rect 392 417788 6188 417816
rect 6244 417788 6254 417844
rect 6402 417676 6412 417732
rect 6468 417676 8120 417732
rect 595560 416836 597000 417032
rect 585554 416780 585564 416836
rect 585620 416808 597000 416836
rect 585620 416780 595672 416808
rect 582008 404236 585452 404292
rect 585508 404236 585518 404292
rect -960 403732 480 403928
rect -960 403704 4172 403732
rect 392 403676 4172 403704
rect 4228 403676 4238 403732
rect 595560 403620 597000 403816
rect 585666 403564 585676 403620
rect 585732 403592 597000 403620
rect 585732 403564 595672 403592
rect 6178 396620 6188 396676
rect 6244 396620 8120 396676
rect 582008 393484 585564 393540
rect 585620 393484 585630 393540
rect 595560 390404 597000 390600
rect 585442 390348 585452 390404
rect 585508 390376 597000 390404
rect 585508 390348 595672 390376
rect -960 389620 480 389816
rect -960 389592 6412 389620
rect 392 389564 6412 389592
rect 6468 389564 6478 389620
rect 4162 386092 4172 386148
rect 4228 386092 8120 386148
rect 582008 382732 585676 382788
rect 585732 382732 585742 382788
rect 595560 377188 597000 377384
rect 585666 377132 585676 377188
rect 585732 377160 597000 377188
rect 585732 377132 595672 377160
rect -960 375508 480 375704
rect 6402 375564 6412 375620
rect 6468 375564 8120 375620
rect -960 375480 6188 375508
rect 392 375452 6188 375480
rect 6244 375452 6254 375508
rect 595560 363972 597000 364168
rect 590482 363916 590492 363972
rect 590548 363944 597000 363972
rect 590548 363916 595672 363944
rect -960 361396 480 361592
rect -960 361368 4172 361396
rect 392 361340 4172 361368
rect 4228 361340 4238 361396
rect 582008 361228 585452 361284
rect 585508 361228 585518 361284
rect 6178 354508 6188 354564
rect 6244 354508 8120 354564
rect 595560 350756 597000 350952
rect 585442 350700 585452 350756
rect 585508 350728 597000 350756
rect 585508 350700 595672 350728
rect 582008 350476 585676 350532
rect 585732 350476 585742 350532
rect -960 347284 480 347480
rect -960 347256 6188 347284
rect 392 347228 6188 347256
rect 6244 347228 6254 347284
rect 4162 343980 4172 344036
rect 4228 343980 8120 344036
rect 582008 339724 590492 339780
rect 590548 339724 590558 339780
rect 595560 337540 597000 337736
rect 585666 337484 585676 337540
rect 585732 337512 597000 337540
rect 585732 337484 595672 337512
rect 6178 333452 6188 333508
rect 6244 333452 8120 333508
rect -960 333172 480 333368
rect -960 333144 4172 333172
rect 392 333116 4172 333144
rect 4228 333116 4238 333172
rect 595560 324324 597000 324520
rect 585554 324268 585564 324324
rect 585620 324296 597000 324324
rect 585620 324268 595672 324296
rect -960 319060 480 319256
rect -960 319032 4284 319060
rect 392 319004 4284 319032
rect 4340 319004 4350 319060
rect 582008 318220 585452 318276
rect 585508 318220 585518 318276
rect 4162 312396 4172 312452
rect 4228 312396 8120 312452
rect 595560 311108 597000 311304
rect 585442 311052 585452 311108
rect 585508 311080 597000 311108
rect 585508 311052 595672 311080
rect 582008 307468 585676 307524
rect 585732 307468 585742 307524
rect -960 304948 480 305144
rect -960 304920 6188 304948
rect 392 304892 6188 304920
rect 6244 304892 6254 304948
rect 4274 301868 4284 301924
rect 4340 301868 8120 301924
rect 595560 297892 597000 298088
rect 590482 297836 590492 297892
rect 590548 297864 597000 297892
rect 590548 297836 595672 297864
rect 582008 296716 585564 296772
rect 585620 296716 585630 296772
rect 6178 291340 6188 291396
rect 6244 291340 8120 291396
rect -960 290836 480 291032
rect -960 290808 4172 290836
rect 392 290780 4172 290808
rect 4228 290780 4238 290836
rect 595560 284676 597000 284872
rect 585554 284620 585564 284676
rect 585620 284648 597000 284676
rect 585620 284620 595672 284648
rect -960 276724 480 276920
rect -960 276696 4284 276724
rect 392 276668 4284 276696
rect 4340 276668 4350 276724
rect 582008 275212 585452 275268
rect 585508 275212 585518 275268
rect 595560 271460 597000 271656
rect 585442 271404 585452 271460
rect 585508 271432 597000 271460
rect 585508 271404 595672 271432
rect 4162 270284 4172 270340
rect 4228 270284 8120 270340
rect 582008 264460 590492 264516
rect 590548 264460 590558 264516
rect -960 262612 480 262808
rect -960 262584 6188 262612
rect 392 262556 6188 262584
rect 6244 262556 6254 262612
rect 4274 259756 4284 259812
rect 4340 259756 8120 259812
rect 595560 258244 597000 258440
rect 587122 258188 587132 258244
rect 587188 258216 597000 258244
rect 587188 258188 595672 258216
rect 582008 253708 585564 253764
rect 585620 253708 585630 253764
rect 6178 249228 6188 249284
rect 6244 249228 8120 249284
rect -960 248500 480 248696
rect -960 248472 6188 248500
rect 392 248444 6188 248472
rect 6244 248444 6254 248500
rect 595560 245028 597000 245224
rect 590482 244972 590492 245028
rect 590548 245000 597000 245028
rect 590548 244972 595672 245000
rect -960 234388 480 234584
rect -960 234360 4172 234388
rect 392 234332 4172 234360
rect 4228 234332 4238 234388
rect 582008 232204 585452 232260
rect 585508 232204 585518 232260
rect 595560 231924 597000 232008
rect 585666 231868 585676 231924
rect 585732 231868 597000 231924
rect 595560 231784 597000 231868
rect 6178 228172 6188 228228
rect 6244 228172 8120 228228
rect 582008 221452 587132 221508
rect 587188 221452 587198 221508
rect -960 220276 480 220472
rect -960 220248 6188 220276
rect 392 220220 6188 220248
rect 6244 220220 6254 220276
rect 595560 218596 597000 218792
rect 585442 218540 585452 218596
rect 585508 218568 597000 218596
rect 585508 218540 595672 218568
rect 4162 217644 4172 217700
rect 4228 217644 8120 217700
rect 582008 210700 590492 210756
rect 590548 210700 590558 210756
rect 6178 207116 6188 207172
rect 6244 207116 8120 207172
rect -960 206164 480 206360
rect -960 206136 6188 206164
rect 392 206108 6188 206136
rect 6244 206108 6254 206164
rect 595560 205380 597000 205576
rect 585554 205324 585564 205380
rect 585620 205352 597000 205380
rect 585620 205324 595672 205352
rect 582008 199948 585676 200004
rect 585732 199948 585742 200004
rect -960 192052 480 192248
rect 595560 192164 597000 192360
rect 585666 192108 585676 192164
rect 585732 192136 597000 192164
rect 585732 192108 595672 192136
rect -960 192024 4172 192052
rect 392 191996 4172 192024
rect 4228 191996 4238 192052
rect 582008 189196 585452 189252
rect 585508 189196 585518 189252
rect 6178 186060 6188 186116
rect 6244 186060 8120 186116
rect 595560 178948 597000 179144
rect 585778 178892 585788 178948
rect 585844 178920 597000 178948
rect 585844 178892 595672 178920
rect 582008 178444 585564 178500
rect 585620 178444 585630 178500
rect -960 177940 480 178136
rect -960 177912 4284 177940
rect 392 177884 4284 177912
rect 4340 177884 4350 177940
rect 4162 175532 4172 175588
rect 4228 175532 8120 175588
rect 582008 167692 585676 167748
rect 585732 167692 585742 167748
rect 595560 165732 597000 165928
rect 585442 165676 585452 165732
rect 585508 165704 597000 165732
rect 585508 165676 595672 165704
rect 4274 165004 4284 165060
rect 4340 165004 8120 165060
rect -960 163828 480 164024
rect -960 163800 6188 163828
rect 392 163772 6188 163800
rect 6244 163772 6254 163828
rect 582008 156940 585788 156996
rect 585844 156940 585854 156996
rect 595560 152516 597000 152712
rect 585554 152460 585564 152516
rect 585620 152488 597000 152516
rect 585620 152460 595672 152488
rect -960 149716 480 149912
rect -960 149688 4172 149716
rect 392 149660 4172 149688
rect 4228 149660 4238 149716
rect 582008 146188 585452 146244
rect 585508 146188 585518 146244
rect 6178 143948 6188 144004
rect 6244 143948 8120 144004
rect 595560 139300 597000 139496
rect 590482 139244 590492 139300
rect 590548 139272 597000 139300
rect 590548 139244 595672 139272
rect -960 135604 480 135800
rect -960 135576 4284 135604
rect 392 135548 4284 135576
rect 4340 135548 4350 135604
rect 582008 135436 585564 135492
rect 585620 135436 585630 135492
rect 4162 133420 4172 133476
rect 4228 133420 8120 133476
rect 595560 126084 597000 126280
rect 590594 126028 590604 126084
rect 590660 126056 597000 126084
rect 590660 126028 595672 126056
rect 582008 124684 590492 124740
rect 590548 124684 590558 124740
rect 4274 122892 4284 122948
rect 4340 122892 8120 122948
rect -960 121492 480 121688
rect -960 121464 4172 121492
rect 392 121436 4172 121464
rect 4228 121436 4238 121492
rect 582008 113932 590604 113988
rect 590660 113932 590670 113988
rect 595560 112868 597000 113064
rect 590818 112812 590828 112868
rect 590884 112840 597000 112868
rect 590884 112812 595672 112840
rect -960 107380 480 107576
rect -960 107352 6188 107380
rect 392 107324 6188 107352
rect 6244 107324 6254 107380
rect 582008 103180 590828 103236
rect 590884 103180 590894 103236
rect 4162 101836 4172 101892
rect 4228 101836 8120 101892
rect 595560 99652 597000 99848
rect 587122 99596 587132 99652
rect 587188 99624 597000 99652
rect 587188 99596 595672 99624
rect -960 93268 480 93464
rect -960 93240 4172 93268
rect 392 93212 4172 93240
rect 4228 93212 4238 93268
rect 582008 92428 587132 92484
rect 587188 92428 587198 92484
rect 6178 91308 6188 91364
rect 6244 91308 8120 91364
rect 595560 86436 597000 86632
rect 590482 86380 590492 86436
rect 590548 86408 597000 86436
rect 590548 86380 595672 86408
rect 582008 81676 590492 81732
rect 590548 81676 590558 81732
rect 4162 80780 4172 80836
rect 4228 80780 8120 80836
rect -960 79156 480 79352
rect -960 79128 4172 79156
rect 392 79100 4172 79128
rect 4228 79100 4238 79156
rect 595560 73220 597000 73416
rect 588914 73164 588924 73220
rect 588980 73192 597000 73220
rect 588980 73164 595672 73192
rect 582008 70924 588924 70980
rect 588980 70924 588990 70980
rect 4162 70252 4172 70308
rect 4228 70252 8120 70308
rect -960 65044 480 65240
rect -960 65016 5068 65044
rect 392 64988 5068 65016
rect 5124 64988 5134 65044
rect 582008 60200 595672 60228
rect 582008 60172 597000 60200
rect 595560 59976 597000 60172
rect 5058 59724 5068 59780
rect 5124 59724 8120 59780
rect -960 50932 480 51128
rect -960 50904 5068 50932
rect 392 50876 5068 50904
rect 5124 50876 5134 50932
rect 582008 49420 590492 49476
rect 590548 49420 590558 49476
rect 5058 49196 5068 49252
rect 5124 49196 8120 49252
rect 590482 46956 590492 47012
rect 590548 46984 595672 47012
rect 590548 46956 597000 46984
rect 595560 46760 597000 46956
rect 4050 38668 4060 38724
rect 4116 38668 8120 38724
rect 582008 38668 588812 38724
rect 588868 38668 588878 38724
rect -960 36932 480 37016
rect -960 36876 4060 36932
rect 4116 36876 4126 36932
rect -960 36792 480 36876
rect 588802 33740 588812 33796
rect 588868 33768 595672 33796
rect 588868 33740 597000 33768
rect 595560 33544 597000 33740
rect 4162 28140 4172 28196
rect 4228 28140 8120 28196
rect 582008 27916 585452 27972
rect 585508 27916 585518 27972
rect 392 22904 4172 22932
rect -960 22876 4172 22904
rect 4228 22876 4238 22932
rect -960 22680 480 22876
rect 595560 20356 597000 20552
rect 585442 20300 585452 20356
rect 585508 20328 597000 20356
rect 585508 20300 595672 20328
rect 6178 17612 6188 17668
rect 6244 17612 8120 17668
rect 582008 17164 585452 17220
rect 585508 17164 585518 17220
rect 392 8792 6188 8820
rect -960 8764 6188 8792
rect 6244 8764 6254 8820
rect -960 8568 480 8764
rect 595560 7140 597000 7336
rect 585442 7084 585452 7140
rect 585508 7112 597000 7140
rect 585508 7084 595672 7112
rect 419458 6636 419468 6692
rect 419524 6636 430332 6692
rect 430388 6636 430398 6692
rect 457090 6636 457100 6692
rect 457156 6636 470204 6692
rect 470260 6636 470270 6692
rect 516226 6636 516236 6692
rect 516292 6636 533036 6692
rect 533092 6636 533102 6692
rect 423042 6524 423052 6580
rect 423108 6524 434028 6580
rect 434084 6524 434094 6580
rect 435586 6524 435596 6580
rect 435652 6524 447356 6580
rect 447412 6524 447422 6580
rect 458882 6524 458892 6580
rect 458948 6524 472108 6580
rect 472164 6524 472174 6580
rect 514434 6524 514444 6580
rect 514500 6524 531132 6580
rect 531188 6524 531198 6580
rect 532354 6524 532364 6580
rect 532420 6524 550172 6580
rect 550228 6524 550238 6580
rect 557414 6524 557452 6580
rect 557508 6524 557518 6580
rect 392578 6412 392588 6468
rect 392644 6412 401660 6468
rect 401716 6412 401726 6468
rect 408706 6412 408716 6468
rect 408772 6412 418796 6468
rect 418852 6412 418862 6468
rect 421250 6412 421260 6468
rect 421316 6412 432124 6468
rect 432180 6412 432190 6468
rect 433794 6412 433804 6468
rect 433860 6412 445452 6468
rect 445508 6412 445518 6468
rect 446338 6412 446348 6468
rect 446404 6412 458780 6468
rect 458836 6412 458846 6468
rect 460674 6412 460684 6468
rect 460740 6412 474012 6468
rect 474068 6412 474078 6468
rect 500098 6412 500108 6468
rect 500164 6412 515900 6468
rect 515956 6412 515966 6468
rect 518018 6412 518028 6468
rect 518084 6412 534940 6468
rect 534996 6412 535006 6468
rect 539522 6412 539532 6468
rect 539588 6412 557788 6468
rect 557844 6412 557854 6468
rect 560998 6412 561036 6468
rect 561092 6412 561102 6468
rect 390786 6300 390796 6356
rect 390852 6300 399868 6356
rect 399924 6300 399944 6356
rect 406914 6300 406924 6356
rect 406980 6300 416892 6356
rect 416948 6300 416958 6356
rect 417666 6300 417676 6356
rect 417732 6300 428428 6356
rect 428484 6300 428494 6356
rect 432002 6300 432012 6356
rect 432068 6300 443548 6356
rect 443604 6300 443614 6356
rect 444546 6300 444556 6356
rect 444612 6300 456988 6356
rect 457044 6300 457054 6356
rect 462466 6300 462476 6356
rect 462532 6300 475916 6356
rect 475972 6300 475982 6356
rect 498306 6300 498316 6356
rect 498372 6300 514108 6356
rect 514164 6300 514174 6356
rect 519810 6300 519820 6356
rect 519876 6300 536844 6356
rect 536900 6300 536910 6356
rect 543106 6300 543116 6356
rect 543172 6300 561596 6356
rect 561652 6300 561662 6356
rect 349570 6188 349580 6244
rect 349636 6188 355964 6244
rect 356020 6188 356030 6244
rect 396162 6188 396172 6244
rect 396228 6188 405468 6244
rect 405524 6188 405534 6244
rect 410498 6188 410508 6244
rect 410564 6188 420700 6244
rect 420756 6188 420766 6244
rect 424834 6188 424844 6244
rect 424900 6188 435932 6244
rect 435988 6188 435998 6244
rect 437378 6188 437388 6244
rect 437444 6188 449260 6244
rect 449316 6188 449326 6244
rect 449922 6188 449932 6244
rect 449988 6188 462588 6244
rect 462644 6188 462654 6244
rect 464258 6188 464268 6244
rect 464324 6188 477820 6244
rect 477876 6188 477886 6244
rect 501890 6188 501900 6244
rect 501956 6188 517804 6244
rect 517860 6188 517870 6244
rect 521602 6188 521612 6244
rect 521668 6188 538748 6244
rect 538804 6188 538814 6244
rect 544898 6188 544908 6244
rect 544964 6188 563500 6244
rect 563556 6188 563566 6244
rect 175298 6076 175308 6132
rect 175364 6076 179340 6132
rect 179396 6076 179406 6132
rect 315522 6076 315532 6132
rect 315588 6076 319788 6132
rect 319844 6076 319854 6132
rect 328066 6076 328076 6132
rect 328132 6076 333116 6132
rect 333172 6076 333182 6132
rect 337026 6076 337036 6132
rect 337092 6076 342748 6132
rect 342804 6076 342814 6132
rect 351362 6076 351372 6132
rect 351428 6076 357868 6132
rect 357924 6076 357934 6132
rect 358530 6076 358540 6132
rect 358596 6076 365484 6132
rect 365540 6076 365550 6132
rect 397954 6076 397964 6132
rect 398020 6076 407372 6132
rect 407428 6076 407438 6132
rect 426626 6076 426636 6132
rect 426692 6076 437836 6132
rect 437892 6076 437902 6132
rect 439170 6076 439180 6132
rect 439236 6076 451164 6132
rect 451220 6076 451230 6132
rect 451714 6076 451724 6132
rect 451780 6076 464492 6132
rect 464548 6076 464558 6132
rect 466050 6076 466060 6132
rect 466116 6076 479724 6132
rect 479780 6076 479790 6132
rect 503682 6076 503692 6132
rect 503748 6076 519708 6132
rect 519764 6076 519774 6132
rect 523394 6076 523404 6132
rect 523460 6076 540652 6132
rect 540708 6076 540718 6132
rect 546690 6076 546700 6132
rect 546756 6076 565404 6132
rect 565460 6076 565470 6132
rect 173394 5964 173404 6020
rect 173460 5964 177548 6020
rect 177604 5964 177614 6020
rect 211474 5964 211484 6020
rect 211540 5964 213388 6020
rect 213444 5964 213454 6020
rect 317314 5964 317324 6020
rect 317380 5964 321692 6020
rect 321748 5964 321758 6020
rect 324482 5964 324492 6020
rect 324548 5964 329308 6020
rect 329364 5964 329384 6020
rect 338818 5964 338828 6020
rect 338884 5964 344540 6020
rect 344596 5964 344606 6020
rect 360322 5964 360332 6020
rect 360388 5964 367388 6020
rect 367444 5964 367454 6020
rect 374658 5964 374668 6020
rect 374724 5964 382620 6020
rect 382676 5964 382686 6020
rect 399746 5964 399756 6020
rect 399812 5964 409276 6020
rect 409332 5964 409342 6020
rect 414082 5964 414092 6020
rect 414148 5964 424508 6020
rect 424564 5964 424574 6020
rect 429090 5964 429100 6020
rect 429156 5964 439740 6020
rect 439796 5964 439806 6020
rect 440962 5964 440972 6020
rect 441028 5964 453068 6020
rect 453124 5964 453134 6020
rect 453506 5964 453516 6020
rect 453572 5964 466396 6020
rect 466452 5964 466462 6020
rect 467842 5964 467852 6020
rect 467908 5964 481628 6020
rect 481684 5964 481694 6020
rect 482178 5964 482188 6020
rect 482244 5964 496860 6020
rect 496916 5964 496926 6020
rect 505474 5964 505484 6020
rect 505540 5964 521612 6020
rect 521668 5964 521678 6020
rect 526978 5964 526988 6020
rect 527044 5964 544460 6020
rect 544516 5964 544526 6020
rect 548482 5964 548492 6020
rect 548548 5964 567308 6020
rect 567364 5964 567374 6020
rect 11554 5852 11564 5908
rect 11620 5852 25228 5908
rect 25284 5852 25294 5908
rect 186722 5852 186732 5908
rect 186788 5852 190092 5908
rect 190148 5852 190158 5908
rect 198146 5852 198156 5908
rect 198212 5852 200844 5908
rect 200900 5852 200910 5908
rect 222898 5852 222908 5908
rect 222964 5852 224140 5908
rect 224196 5852 224206 5908
rect 258178 5852 258188 5908
rect 258244 5852 258860 5908
rect 258916 5852 258926 5908
rect 281474 5852 281484 5908
rect 281540 5852 283612 5908
rect 283668 5852 283678 5908
rect 313730 5852 313740 5908
rect 313796 5852 317884 5908
rect 317940 5852 317950 5908
rect 326274 5852 326284 5908
rect 326340 5852 331212 5908
rect 331268 5852 331278 5908
rect 340610 5852 340620 5908
rect 340676 5852 346444 5908
rect 346500 5852 346510 5908
rect 347778 5852 347788 5908
rect 347844 5852 354060 5908
rect 354116 5852 354126 5908
rect 362114 5852 362124 5908
rect 362180 5852 369292 5908
rect 369348 5852 369358 5908
rect 394370 5852 394380 5908
rect 394436 5852 403564 5908
rect 403620 5852 403630 5908
rect 405122 5852 405132 5908
rect 405188 5852 414988 5908
rect 415044 5852 415054 5908
rect 415874 5852 415884 5908
rect 415940 5852 426412 5908
rect 426468 5852 426478 5908
rect 430210 5852 430220 5908
rect 430276 5852 441644 5908
rect 441700 5852 441710 5908
rect 442754 5852 442764 5908
rect 442820 5852 454972 5908
rect 455028 5852 455038 5908
rect 455298 5852 455308 5908
rect 455364 5852 468300 5908
rect 468356 5852 468366 5908
rect 469634 5852 469644 5908
rect 469700 5852 483532 5908
rect 483588 5852 483598 5908
rect 483970 5852 483980 5908
rect 484036 5852 498764 5908
rect 498820 5852 498830 5908
rect 507266 5852 507276 5908
rect 507332 5852 523516 5908
rect 523572 5852 523582 5908
rect 528770 5852 528780 5908
rect 528836 5852 546364 5908
rect 546420 5852 546430 5908
rect 550274 5852 550284 5908
rect 550340 5852 569212 5908
rect 569268 5852 569278 5908
rect 448130 5740 448140 5796
rect 448196 5740 460684 5796
rect 460740 5740 460750 5796
rect 512642 5740 512652 5796
rect 512708 5740 529228 5796
rect 529284 5740 529294 5796
rect 277890 5404 277900 5460
rect 277956 5404 279804 5460
rect 279860 5404 279870 5460
rect 177202 5292 177212 5348
rect 177268 5292 181132 5348
rect 181188 5292 181198 5348
rect 333442 5292 333452 5348
rect 333508 5292 338828 5348
rect 338884 5292 338894 5348
rect 345986 5292 345996 5348
rect 346052 5292 352156 5348
rect 352212 5292 352222 5348
rect 356738 5292 356748 5348
rect 356804 5292 363580 5348
rect 363636 5292 363646 5348
rect 179106 5180 179116 5236
rect 179172 5180 182924 5236
rect 182980 5180 182990 5236
rect 190530 5180 190540 5236
rect 190596 5180 193676 5236
rect 193732 5180 193742 5236
rect 194338 5180 194348 5236
rect 194404 5180 197260 5236
rect 197316 5180 197326 5236
rect 200050 5180 200060 5236
rect 200116 5180 202636 5236
rect 202692 5180 202702 5236
rect 203858 5180 203868 5236
rect 203924 5180 206220 5236
rect 206276 5180 206286 5236
rect 207666 5180 207676 5236
rect 207732 5180 209804 5236
rect 209860 5180 209870 5236
rect 213266 5180 213276 5236
rect 213332 5180 215180 5236
rect 215236 5180 215246 5236
rect 276098 5180 276108 5236
rect 276164 5180 277900 5236
rect 277956 5180 277966 5236
rect 295810 5180 295820 5236
rect 295876 5180 298844 5236
rect 298900 5180 298910 5236
rect 311938 5180 311948 5236
rect 312004 5180 315980 5236
rect 316036 5180 316046 5236
rect 331650 5180 331660 5236
rect 331716 5180 336924 5236
rect 336980 5180 336990 5236
rect 344194 5180 344204 5236
rect 344260 5180 350252 5236
rect 350308 5180 350318 5236
rect 354946 5180 354956 5236
rect 355012 5180 361676 5236
rect 361732 5180 361742 5236
rect 171490 5068 171500 5124
rect 171556 5068 175756 5124
rect 175812 5068 175822 5124
rect 181010 5068 181020 5124
rect 181076 5068 184716 5124
rect 184772 5068 184782 5124
rect 188626 5068 188636 5124
rect 188692 5068 191884 5124
rect 191940 5068 191950 5124
rect 192434 5068 192444 5124
rect 192500 5068 195468 5124
rect 195524 5068 195534 5124
rect 196242 5068 196252 5124
rect 196308 5068 199052 5124
rect 199108 5068 199118 5124
rect 201954 5068 201964 5124
rect 202020 5068 204428 5124
rect 204484 5068 204494 5124
rect 205762 5068 205772 5124
rect 205828 5068 208012 5124
rect 208068 5068 208078 5124
rect 209570 5068 209580 5124
rect 209636 5068 211596 5124
rect 211652 5068 211662 5124
rect 215282 5068 215292 5124
rect 215348 5068 216972 5124
rect 217028 5068 217038 5124
rect 217186 5068 217196 5124
rect 217252 5068 218764 5124
rect 218820 5068 218830 5124
rect 265346 5068 265356 5124
rect 265412 5068 266476 5124
rect 266532 5068 266542 5124
rect 270722 5068 270732 5124
rect 270788 5068 272188 5124
rect 272244 5068 272254 5124
rect 272514 5068 272524 5124
rect 272580 5068 274092 5124
rect 274148 5068 274158 5124
rect 274306 5068 274316 5124
rect 274372 5068 275996 5124
rect 276052 5068 276062 5124
rect 279682 5068 279692 5124
rect 279748 5068 281708 5124
rect 281764 5068 281774 5124
rect 294018 5068 294028 5124
rect 294084 5068 296940 5124
rect 296996 5068 297006 5124
rect 310146 5068 310156 5124
rect 310212 5068 314188 5124
rect 314244 5068 314254 5124
rect 319106 5068 319116 5124
rect 319172 5068 323596 5124
rect 323652 5068 323662 5124
rect 329858 5068 329868 5124
rect 329924 5068 335020 5124
rect 335076 5068 335086 5124
rect 335234 5068 335244 5124
rect 335300 5068 340732 5124
rect 340788 5068 340798 5124
rect 342402 5068 342412 5124
rect 342468 5068 348348 5124
rect 348404 5068 348414 5124
rect 353154 5068 353164 5124
rect 353220 5068 359772 5124
rect 359828 5068 359838 5124
rect 376450 5068 376460 5124
rect 376516 5068 384524 5124
rect 384580 5068 384590 5124
rect 412290 5068 412300 5124
rect 412356 5068 422604 5124
rect 422660 5068 422670 5124
rect 26786 4956 26796 5012
rect 26852 4956 39564 5012
rect 39620 4956 39630 5012
rect 64866 4956 64876 5012
rect 64932 4956 75404 5012
rect 75460 4956 75470 5012
rect 24882 4844 24892 4900
rect 24948 4844 37772 4900
rect 37828 4844 37838 4900
rect 41906 4844 41916 4900
rect 41972 4844 53900 4900
rect 53956 4844 53966 4900
rect 55346 4844 55356 4900
rect 55412 4844 66444 4900
rect 66500 4844 66510 4900
rect 485762 4844 485772 4900
rect 485828 4844 500668 4900
rect 500724 4844 500734 4900
rect 534146 4844 534156 4900
rect 534212 4844 552188 4900
rect 552244 4844 552254 4900
rect 22978 4732 22988 4788
rect 23044 4732 35980 4788
rect 36036 4732 36046 4788
rect 40114 4732 40124 4788
rect 40180 4732 52108 4788
rect 52164 4732 52174 4788
rect 53442 4732 53452 4788
rect 53508 4732 64652 4788
rect 64708 4732 64718 4788
rect 76290 4732 76300 4788
rect 76356 4732 86156 4788
rect 86212 4732 86222 4788
rect 87714 4732 87724 4788
rect 87780 4732 96908 4788
rect 96964 4732 96974 4788
rect 125794 4732 125804 4788
rect 125860 4732 132748 4788
rect 132804 4732 132814 4788
rect 473218 4732 473228 4788
rect 473284 4732 487340 4788
rect 487396 4732 487406 4788
rect 487554 4732 487564 4788
rect 487620 4732 502572 4788
rect 502628 4732 502638 4788
rect 553858 4732 553868 4788
rect 553924 4732 573020 4788
rect 573076 4732 573086 4788
rect 21074 4620 21084 4676
rect 21140 4620 34188 4676
rect 34244 4620 34254 4676
rect 38210 4620 38220 4676
rect 38276 4620 50316 4676
rect 50372 4620 50382 4676
rect 51538 4620 51548 4676
rect 51604 4620 62860 4676
rect 62916 4620 62926 4676
rect 66770 4620 66780 4676
rect 66836 4620 77196 4676
rect 77252 4620 77262 4676
rect 78194 4620 78204 4676
rect 78260 4620 87948 4676
rect 88004 4620 88014 4676
rect 89618 4620 89628 4676
rect 89684 4620 98700 4676
rect 98756 4620 98766 4676
rect 104850 4620 104860 4676
rect 104916 4620 113036 4676
rect 113092 4620 113102 4676
rect 114370 4620 114380 4676
rect 114436 4620 121996 4676
rect 122052 4620 122062 4676
rect 123890 4620 123900 4676
rect 123956 4620 130956 4676
rect 131012 4620 131022 4676
rect 146738 4620 146748 4676
rect 146804 4620 152460 4676
rect 152516 4620 152526 4676
rect 308354 4620 308364 4676
rect 308420 4620 312172 4676
rect 312228 4620 312238 4676
rect 381826 4620 381836 4676
rect 381892 4620 390236 4676
rect 390292 4620 390302 4676
rect 471426 4620 471436 4676
rect 471492 4620 485548 4676
rect 485604 4620 485614 4676
rect 489346 4620 489356 4676
rect 489412 4620 504476 4676
rect 504532 4620 504542 4676
rect 525186 4620 525196 4676
rect 525252 4620 542668 4676
rect 542724 4620 542734 4676
rect 552066 4620 552076 4676
rect 552132 4620 571228 4676
rect 571284 4620 571294 4676
rect 19170 4508 19180 4564
rect 19236 4508 32396 4564
rect 32452 4508 32462 4564
rect 36306 4508 36316 4564
rect 36372 4508 48524 4564
rect 48580 4508 48590 4564
rect 49634 4508 49644 4564
rect 49700 4508 61068 4564
rect 61124 4508 61134 4564
rect 62962 4508 62972 4564
rect 63028 4508 73612 4564
rect 73668 4508 73678 4564
rect 74386 4508 74396 4564
rect 74452 4508 84364 4564
rect 84420 4508 84430 4564
rect 85810 4508 85820 4564
rect 85876 4508 95116 4564
rect 95172 4508 95182 4564
rect 99026 4508 99036 4564
rect 99092 4508 107660 4564
rect 107716 4508 107726 4564
rect 141026 4508 141036 4564
rect 141092 4508 147084 4564
rect 147140 4508 147150 4564
rect 148642 4508 148652 4564
rect 148708 4508 154252 4564
rect 154308 4508 154318 4564
rect 383618 4508 383628 4564
rect 383684 4508 392140 4564
rect 392196 4508 392206 4564
rect 475010 4508 475020 4564
rect 475076 4508 489244 4564
rect 489300 4508 489310 4564
rect 491138 4508 491148 4564
rect 491204 4508 506380 4564
rect 506436 4508 506446 4564
rect 530562 4508 530572 4564
rect 530628 4508 548268 4564
rect 548324 4508 548334 4564
rect 555650 4508 555660 4564
rect 555716 4508 574924 4564
rect 574980 4508 574990 4564
rect 17266 4396 17276 4452
rect 17332 4396 30604 4452
rect 30660 4396 30670 4452
rect 34402 4396 34412 4452
rect 34468 4396 46732 4452
rect 46788 4396 46798 4452
rect 47730 4396 47740 4452
rect 47796 4396 59276 4452
rect 59332 4396 59342 4452
rect 61170 4396 61180 4452
rect 61236 4396 71820 4452
rect 71876 4396 71886 4452
rect 72482 4396 72492 4452
rect 72548 4396 82572 4452
rect 82628 4396 82638 4452
rect 97234 4396 97244 4452
rect 97300 4396 105868 4452
rect 105924 4396 105934 4452
rect 116274 4396 116284 4452
rect 116340 4396 123788 4452
rect 123844 4396 123854 4452
rect 127586 4396 127596 4452
rect 127652 4396 134540 4452
rect 134596 4396 134606 4452
rect 135314 4396 135324 4452
rect 135380 4396 141708 4452
rect 141764 4396 141774 4452
rect 150546 4396 150556 4452
rect 150612 4396 156044 4452
rect 156100 4396 156110 4452
rect 163874 4396 163884 4452
rect 163940 4396 168588 4452
rect 168644 4396 168654 4452
rect 304770 4396 304780 4452
rect 304836 4396 308364 4452
rect 308420 4396 308430 4452
rect 363906 4396 363916 4452
rect 363972 4396 371308 4452
rect 371364 4396 371374 4452
rect 372866 4396 372876 4452
rect 372932 4396 380716 4452
rect 380772 4396 380782 4452
rect 385410 4396 385420 4452
rect 385476 4396 394044 4452
rect 394100 4396 394110 4452
rect 480386 4396 480396 4452
rect 480452 4396 494956 4452
rect 495012 4396 495022 4452
rect 496514 4396 496524 4452
rect 496580 4396 512092 4452
rect 512148 4396 512158 4452
rect 535938 4396 535948 4452
rect 536004 4396 553980 4452
rect 554036 4396 554046 4452
rect 562818 4396 562828 4452
rect 562884 4396 582540 4452
rect 582596 4396 582606 4452
rect 15362 4284 15372 4340
rect 15428 4284 28812 4340
rect 28868 4284 28878 4340
rect 32498 4284 32508 4340
rect 32564 4284 44940 4340
rect 44996 4284 45006 4340
rect 45826 4284 45836 4340
rect 45892 4284 57484 4340
rect 57540 4284 57550 4340
rect 70466 4284 70476 4340
rect 70532 4284 80780 4340
rect 80836 4284 80846 4340
rect 82002 4284 82012 4340
rect 82068 4284 90860 4340
rect 90916 4284 90926 4340
rect 93426 4284 93436 4340
rect 93492 4284 102284 4340
rect 102340 4284 102350 4340
rect 102946 4284 102956 4340
rect 103012 4284 111244 4340
rect 111300 4284 111310 4340
rect 112466 4284 112476 4340
rect 112532 4284 120204 4340
rect 120260 4284 120270 4340
rect 139122 4284 139132 4340
rect 139188 4284 145292 4340
rect 145348 4284 145358 4340
rect 161970 4284 161980 4340
rect 162036 4284 166796 4340
rect 166852 4284 166862 4340
rect 184706 4284 184716 4340
rect 184772 4284 188300 4340
rect 188356 4284 188366 4340
rect 369506 4284 369516 4340
rect 369572 4284 376908 4340
rect 376964 4284 376974 4340
rect 387202 4284 387212 4340
rect 387268 4284 395948 4340
rect 396004 4284 396014 4340
rect 476802 4284 476812 4340
rect 476868 4284 491148 4340
rect 491204 4284 491214 4340
rect 492930 4284 492940 4340
rect 492996 4284 508284 4340
rect 508340 4284 508350 4340
rect 509058 4284 509068 4340
rect 509124 4284 525420 4340
rect 525476 4284 525486 4340
rect 541314 4284 541324 4340
rect 541380 4284 559692 4340
rect 559748 4284 559758 4340
rect 564610 4284 564620 4340
rect 564676 4284 584444 4340
rect 584500 4284 584510 4340
rect 13346 4172 13356 4228
rect 13412 4172 27020 4228
rect 27076 4172 27086 4228
rect 30594 4172 30604 4228
rect 30660 4172 43148 4228
rect 43204 4172 43214 4228
rect 43922 4172 43932 4228
rect 43988 4172 55692 4228
rect 55748 4172 55758 4228
rect 57250 4172 57260 4228
rect 57316 4172 68236 4228
rect 68292 4172 68302 4228
rect 68674 4172 68684 4228
rect 68740 4172 78988 4228
rect 79044 4172 79054 4228
rect 80098 4172 80108 4228
rect 80164 4172 89740 4228
rect 89796 4172 89806 4228
rect 91522 4172 91532 4228
rect 91588 4172 100492 4228
rect 100548 4172 100558 4228
rect 101042 4172 101052 4228
rect 101108 4172 109452 4228
rect 109508 4172 109518 4228
rect 110562 4172 110572 4228
rect 110628 4172 118412 4228
rect 118468 4172 118478 4228
rect 129602 4172 129612 4228
rect 129668 4172 136332 4228
rect 136388 4172 136398 4228
rect 137218 4172 137228 4228
rect 137284 4172 143500 4228
rect 143556 4172 143566 4228
rect 152450 4172 152460 4228
rect 152516 4172 157836 4228
rect 157892 4172 157902 4228
rect 160066 4172 160076 4228
rect 160132 4172 165004 4228
rect 165060 4172 165070 4228
rect 165778 4172 165788 4228
rect 165844 4172 170380 4228
rect 170436 4172 170446 4228
rect 292226 4172 292236 4228
rect 292292 4172 295036 4228
rect 295092 4172 295102 4228
rect 302978 4172 302988 4228
rect 303044 4172 306460 4228
rect 306516 4172 306526 4228
rect 371074 4172 371084 4228
rect 371140 4172 378812 4228
rect 378868 4172 378878 4228
rect 380034 4172 380044 4228
rect 380100 4172 388332 4228
rect 388388 4172 388398 4228
rect 403330 4172 403340 4228
rect 403396 4172 413084 4228
rect 413140 4172 413150 4228
rect 478594 4172 478604 4228
rect 478660 4172 493052 4228
rect 493108 4172 493118 4228
rect 494722 4172 494732 4228
rect 494788 4172 510188 4228
rect 510244 4172 510254 4228
rect 510850 4172 510860 4228
rect 510916 4172 527324 4228
rect 527380 4172 527390 4228
rect 537730 4172 537740 4228
rect 537796 4172 555884 4228
rect 555940 4172 555950 4228
rect 559234 4172 559244 4228
rect 559300 4172 578732 4228
rect 578788 4172 578798 4228
rect 28690 4060 28700 4116
rect 28756 4060 41356 4116
rect 41412 4060 41422 4116
rect 59154 4060 59164 4116
rect 59220 4060 70028 4116
rect 70084 4060 70094 4116
rect 83906 4060 83916 4116
rect 83972 4060 93324 4116
rect 93380 4060 93390 4116
rect 95330 4060 95340 4116
rect 95396 4060 104076 4116
rect 104132 4060 104142 4116
rect 108658 4060 108668 4116
rect 108724 4060 116620 4116
rect 116676 4060 116686 4116
rect 121986 4060 121996 4116
rect 122052 4060 129164 4116
rect 129220 4060 129230 4116
rect 133410 4060 133420 4116
rect 133476 4060 139916 4116
rect 139972 4060 139982 4116
rect 144834 4060 144844 4116
rect 144900 4060 150668 4116
rect 150724 4060 150734 4116
rect 158162 4060 158172 4116
rect 158228 4060 163212 4116
rect 163268 4060 163278 4116
rect 169586 4060 169596 4116
rect 169652 4060 173964 4116
rect 174020 4060 174030 4116
rect 182914 4060 182924 4116
rect 182980 4060 186508 4116
rect 186564 4060 186574 4116
rect 283266 4060 283276 4116
rect 283332 4060 285628 4116
rect 285684 4060 285694 4116
rect 286850 4060 286860 4116
rect 286916 4060 289324 4116
rect 289380 4060 289390 4116
rect 290434 4060 290444 4116
rect 290500 4060 293132 4116
rect 293188 4060 293198 4116
rect 297602 4060 297612 4116
rect 297668 4060 300748 4116
rect 300804 4060 300814 4116
rect 301186 4060 301196 4116
rect 301252 4060 304556 4116
rect 304612 4060 304622 4116
rect 306562 4060 306572 4116
rect 306628 4060 310268 4116
rect 310324 4060 310334 4116
rect 320898 4060 320908 4116
rect 320964 4060 325500 4116
rect 325556 4060 325566 4116
rect 365698 4060 365708 4116
rect 365764 4060 373100 4116
rect 373156 4060 373166 4116
rect 378242 4060 378252 4116
rect 378308 4060 386428 4116
rect 386484 4060 386494 4116
rect 388994 4060 389004 4116
rect 389060 4060 397852 4116
rect 397908 4060 397918 4116
rect 401538 4060 401548 4116
rect 401604 4060 411180 4116
rect 411236 4060 411246 4116
rect 106754 3948 106764 4004
rect 106820 3948 114828 4004
rect 114884 3948 114894 4004
rect 120082 3948 120092 4004
rect 120148 3948 127372 4004
rect 127428 3948 127438 4004
rect 131506 3948 131516 4004
rect 131572 3948 138124 4004
rect 138180 3948 138190 4004
rect 142930 3948 142940 4004
rect 142996 3948 148876 4004
rect 148932 3948 148942 4004
rect 156146 3948 156156 4004
rect 156212 3948 161420 4004
rect 161476 3948 161486 4004
rect 167682 3948 167692 4004
rect 167748 3948 172172 4004
rect 172228 3948 172238 4004
rect 285058 3948 285068 4004
rect 285124 3948 287420 4004
rect 287476 3948 287486 4004
rect 288642 3948 288652 4004
rect 288708 3948 291228 4004
rect 291284 3948 291294 4004
rect 299394 3948 299404 4004
rect 299460 3948 302652 4004
rect 302708 3948 302718 4004
rect 322690 3948 322700 4004
rect 322756 3948 327404 4004
rect 327460 3948 327470 4004
rect 367490 3948 367500 4004
rect 367556 3948 375004 4004
rect 375060 3948 375070 4004
rect 118178 3836 118188 3892
rect 118244 3836 125580 3892
rect 125636 3836 125646 3892
rect 154354 3836 154364 3892
rect 154420 3836 159628 3892
rect 159684 3836 159694 3892
rect 576790 3388 576828 3444
rect 576884 3388 576894 3444
rect 580598 3388 580636 3444
rect 580692 3388 580702 3444
<< via3 >>
rect 590492 588588 590548 588644
rect 4172 587132 4228 587188
rect 590492 576268 590548 576324
rect 591276 575372 591332 575428
rect 4284 573020 4340 573076
rect 591276 565516 591332 565572
rect 4172 565068 4228 565124
rect 586348 562156 586404 562212
rect 6188 558908 6244 558964
rect 586348 554764 586404 554820
rect 4284 554540 4340 554596
rect 590492 548940 590548 548996
rect 4172 544796 4228 544852
rect 6188 544012 6244 544068
rect 588588 535724 588644 535780
rect 590492 533260 590548 533316
rect 4284 530684 4340 530740
rect 4172 522956 4228 523012
rect 588588 522508 588644 522564
rect 588812 522508 588868 522564
rect 6188 516572 6244 516628
rect 4284 512428 4340 512484
rect 588812 511756 588868 511812
rect 585452 509292 585508 509348
rect 4172 502460 4228 502516
rect 6188 501900 6244 501956
rect 590492 496076 590548 496132
rect 585452 490252 585508 490308
rect 4284 488348 4340 488404
rect 590604 482860 590660 482916
rect 4172 480844 4228 480900
rect 590492 479500 590548 479556
rect 6412 474236 6468 474292
rect 4284 470316 4340 470372
rect 585452 469644 585508 469700
rect 590604 468748 590660 468804
rect 6188 460124 6244 460180
rect 6412 459788 6468 459844
rect 585564 456428 585620 456484
rect 585452 447244 585508 447300
rect 4172 446012 4228 446068
rect 590492 443212 590548 443268
rect 6188 438732 6244 438788
rect 585564 436492 585620 436548
rect 6412 431900 6468 431956
rect 585452 430108 585508 430164
rect 4172 428204 4228 428260
rect 590492 425740 590548 425796
rect 6188 417788 6244 417844
rect 6412 417676 6468 417732
rect 585564 416780 585620 416836
rect 585452 404236 585508 404292
rect 4172 403676 4228 403732
rect 585676 403564 585732 403620
rect 6188 396620 6244 396676
rect 585564 393484 585620 393540
rect 585452 390348 585508 390404
rect 6412 389564 6468 389620
rect 4172 386092 4228 386148
rect 585676 382732 585732 382788
rect 585676 377132 585732 377188
rect 6412 375564 6468 375620
rect 6188 375452 6244 375508
rect 590492 363916 590548 363972
rect 4172 361340 4228 361396
rect 585452 361228 585508 361284
rect 6188 354508 6244 354564
rect 585452 350700 585508 350756
rect 585676 350476 585732 350532
rect 6188 347228 6244 347284
rect 4172 343980 4228 344036
rect 590492 339724 590548 339780
rect 585676 337484 585732 337540
rect 6188 333452 6244 333508
rect 4172 333116 4228 333172
rect 585564 324268 585620 324324
rect 4284 319004 4340 319060
rect 585452 318220 585508 318276
rect 4172 312396 4228 312452
rect 585452 311052 585508 311108
rect 585676 307468 585732 307524
rect 6188 304892 6244 304948
rect 4284 301868 4340 301924
rect 590492 297836 590548 297892
rect 585564 296716 585620 296772
rect 6188 291340 6244 291396
rect 4172 290780 4228 290836
rect 585564 284620 585620 284676
rect 4284 276668 4340 276724
rect 585452 275212 585508 275268
rect 585452 271404 585508 271460
rect 4172 270284 4228 270340
rect 590492 264460 590548 264516
rect 6188 262556 6244 262612
rect 4284 259756 4340 259812
rect 587132 258188 587188 258244
rect 585564 253708 585620 253764
rect 6188 249228 6244 249284
rect 6188 248444 6244 248500
rect 590492 244972 590548 245028
rect 4172 234332 4228 234388
rect 585452 232204 585508 232260
rect 585676 231868 585732 231924
rect 6188 228172 6244 228228
rect 587132 221452 587188 221508
rect 6188 220220 6244 220276
rect 585452 218540 585508 218596
rect 4172 217644 4228 217700
rect 590492 210700 590548 210756
rect 6188 207116 6244 207172
rect 6188 206108 6244 206164
rect 585564 205324 585620 205380
rect 585676 199948 585732 200004
rect 585676 192108 585732 192164
rect 4172 191996 4228 192052
rect 585452 189196 585508 189252
rect 6188 186060 6244 186116
rect 585788 178892 585844 178948
rect 585564 178444 585620 178500
rect 4284 177884 4340 177940
rect 4172 175532 4228 175588
rect 585676 167692 585732 167748
rect 585452 165676 585508 165732
rect 4284 165004 4340 165060
rect 6188 163772 6244 163828
rect 585788 156940 585844 156996
rect 585564 152460 585620 152516
rect 4172 149660 4228 149716
rect 585452 146188 585508 146244
rect 6188 143948 6244 144004
rect 590492 139244 590548 139300
rect 4284 135548 4340 135604
rect 585564 135436 585620 135492
rect 4172 133420 4228 133476
rect 590604 126028 590660 126084
rect 590492 124684 590548 124740
rect 4284 122892 4340 122948
rect 4172 121436 4228 121492
rect 590604 113932 590660 113988
rect 590828 112812 590884 112868
rect 6188 107324 6244 107380
rect 590828 103180 590884 103236
rect 4172 101836 4228 101892
rect 587132 99596 587188 99652
rect 4172 93212 4228 93268
rect 587132 92428 587188 92484
rect 6188 91308 6244 91364
rect 590492 86380 590548 86436
rect 590492 81676 590548 81732
rect 4172 80780 4228 80836
rect 4172 79100 4228 79156
rect 588924 73164 588980 73220
rect 588924 70924 588980 70980
rect 4172 70252 4228 70308
rect 5068 64988 5124 65044
rect 5068 59724 5124 59780
rect 5068 50876 5124 50932
rect 590492 49420 590548 49476
rect 5068 49196 5124 49252
rect 590492 46956 590548 47012
rect 4060 38668 4116 38724
rect 588812 38668 588868 38724
rect 4060 36876 4116 36932
rect 588812 33740 588868 33796
rect 4172 28140 4228 28196
rect 585452 27916 585508 27972
rect 4172 22876 4228 22932
rect 585452 20300 585508 20356
rect 6188 17612 6244 17668
rect 585452 17164 585508 17220
rect 6188 8764 6244 8820
rect 585452 7084 585508 7140
rect 557452 6524 557508 6580
rect 561036 6412 561092 6468
rect 576828 3388 576884 3444
rect 580636 3388 580692 3444
<< metal4 >>
rect -1916 598172 -1296 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 -1296 598172
rect -1916 598048 -1296 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 -1296 598048
rect -1916 597924 -1296 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 -1296 597924
rect -1916 597800 -1296 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 -1296 597800
rect -1916 586350 -1296 597744
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 -1296 586350
rect -1916 586226 -1296 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 -1296 586226
rect -1916 586102 -1296 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 -1296 586102
rect -1916 585978 -1296 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 -1296 585978
rect -1916 568350 -1296 585922
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 -1296 568350
rect -1916 568226 -1296 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 -1296 568226
rect -1916 568102 -1296 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 -1296 568102
rect -1916 567978 -1296 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 -1296 567978
rect -1916 550350 -1296 567922
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 -1296 550350
rect -1916 550226 -1296 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 -1296 550226
rect -1916 550102 -1296 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 -1296 550102
rect -1916 549978 -1296 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 -1296 549978
rect -1916 532350 -1296 549922
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 -1296 532350
rect -1916 532226 -1296 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 -1296 532226
rect -1916 532102 -1296 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 -1296 532102
rect -1916 531978 -1296 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 -1296 531978
rect -1916 514350 -1296 531922
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 -1296 514350
rect -1916 514226 -1296 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 -1296 514226
rect -1916 514102 -1296 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 -1296 514102
rect -1916 513978 -1296 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 -1296 513978
rect -1916 496350 -1296 513922
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 -1296 496350
rect -1916 496226 -1296 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 -1296 496226
rect -1916 496102 -1296 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 -1296 496102
rect -1916 495978 -1296 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 -1296 495978
rect -1916 478350 -1296 495922
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 -1296 478350
rect -1916 478226 -1296 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 -1296 478226
rect -1916 478102 -1296 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 -1296 478102
rect -1916 477978 -1296 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 -1296 477978
rect -1916 460350 -1296 477922
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 -1296 460350
rect -1916 460226 -1296 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 -1296 460226
rect -1916 460102 -1296 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 -1296 460102
rect -1916 459978 -1296 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 -1296 459978
rect -1916 442350 -1296 459922
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 -1296 442350
rect -1916 442226 -1296 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 -1296 442226
rect -1916 442102 -1296 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 -1296 442102
rect -1916 441978 -1296 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 -1296 441978
rect -1916 424350 -1296 441922
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 -1296 424350
rect -1916 424226 -1296 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 -1296 424226
rect -1916 424102 -1296 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 -1296 424102
rect -1916 423978 -1296 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 -1296 423978
rect -1916 406350 -1296 423922
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 -1296 406350
rect -1916 406226 -1296 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 -1296 406226
rect -1916 406102 -1296 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 -1296 406102
rect -1916 405978 -1296 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 -1296 405978
rect -1916 388350 -1296 405922
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 -1296 388350
rect -1916 388226 -1296 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 -1296 388226
rect -1916 388102 -1296 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 -1296 388102
rect -1916 387978 -1296 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 -1296 387978
rect -1916 370350 -1296 387922
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 -1296 370350
rect -1916 370226 -1296 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 -1296 370226
rect -1916 370102 -1296 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 -1296 370102
rect -1916 369978 -1296 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 -1296 369978
rect -1916 352350 -1296 369922
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 -1296 352350
rect -1916 352226 -1296 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 -1296 352226
rect -1916 352102 -1296 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 -1296 352102
rect -1916 351978 -1296 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 -1296 351978
rect -1916 334350 -1296 351922
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 -1296 334350
rect -1916 334226 -1296 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 -1296 334226
rect -1916 334102 -1296 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 -1296 334102
rect -1916 333978 -1296 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 -1296 333978
rect -1916 316350 -1296 333922
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 -1296 316350
rect -1916 316226 -1296 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 -1296 316226
rect -1916 316102 -1296 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 -1296 316102
rect -1916 315978 -1296 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 -1296 315978
rect -1916 298350 -1296 315922
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 -1296 298350
rect -1916 298226 -1296 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 -1296 298226
rect -1916 298102 -1296 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 -1296 298102
rect -1916 297978 -1296 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 -1296 297978
rect -1916 280350 -1296 297922
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 -1296 280350
rect -1916 280226 -1296 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 -1296 280226
rect -1916 280102 -1296 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 -1296 280102
rect -1916 279978 -1296 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 -1296 279978
rect -1916 262350 -1296 279922
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 -1296 262350
rect -1916 262226 -1296 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 -1296 262226
rect -1916 262102 -1296 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 -1296 262102
rect -1916 261978 -1296 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 -1296 261978
rect -1916 244350 -1296 261922
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 -1296 244350
rect -1916 244226 -1296 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 -1296 244226
rect -1916 244102 -1296 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 -1296 244102
rect -1916 243978 -1296 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 -1296 243978
rect -1916 226350 -1296 243922
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 -1296 226350
rect -1916 226226 -1296 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 -1296 226226
rect -1916 226102 -1296 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 -1296 226102
rect -1916 225978 -1296 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 -1296 225978
rect -1916 208350 -1296 225922
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 -1296 208350
rect -1916 208226 -1296 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 -1296 208226
rect -1916 208102 -1296 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 -1296 208102
rect -1916 207978 -1296 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 -1296 207978
rect -1916 190350 -1296 207922
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 -1296 190350
rect -1916 190226 -1296 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 -1296 190226
rect -1916 190102 -1296 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 -1296 190102
rect -1916 189978 -1296 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 -1296 189978
rect -1916 172350 -1296 189922
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 -1296 172350
rect -1916 172226 -1296 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 -1296 172226
rect -1916 172102 -1296 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 -1296 172102
rect -1916 171978 -1296 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 -1296 171978
rect -1916 154350 -1296 171922
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 -1296 154350
rect -1916 154226 -1296 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 -1296 154226
rect -1916 154102 -1296 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 -1296 154102
rect -1916 153978 -1296 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 -1296 153978
rect -1916 136350 -1296 153922
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 -1296 136350
rect -1916 136226 -1296 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 -1296 136226
rect -1916 136102 -1296 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 -1296 136102
rect -1916 135978 -1296 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 -1296 135978
rect -1916 118350 -1296 135922
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 -1296 118350
rect -1916 118226 -1296 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 -1296 118226
rect -1916 118102 -1296 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 -1296 118102
rect -1916 117978 -1296 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 -1296 117978
rect -1916 100350 -1296 117922
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 -1296 100350
rect -1916 100226 -1296 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 -1296 100226
rect -1916 100102 -1296 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 -1296 100102
rect -1916 99978 -1296 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 -1296 99978
rect -1916 82350 -1296 99922
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 -1296 82350
rect -1916 82226 -1296 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 -1296 82226
rect -1916 82102 -1296 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 -1296 82102
rect -1916 81978 -1296 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 -1296 81978
rect -1916 64350 -1296 81922
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 -1296 64350
rect -1916 64226 -1296 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 -1296 64226
rect -1916 64102 -1296 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 -1296 64102
rect -1916 63978 -1296 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 -1296 63978
rect -1916 46350 -1296 63922
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 -1296 46350
rect -1916 46226 -1296 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 -1296 46226
rect -1916 46102 -1296 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 -1296 46102
rect -1916 45978 -1296 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 -1296 45978
rect -1916 28350 -1296 45922
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 -1296 28350
rect -1916 28226 -1296 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 -1296 28226
rect -1916 28102 -1296 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 -1296 28102
rect -1916 27978 -1296 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 -1296 27978
rect -1916 10350 -1296 27922
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 -1296 10350
rect -1916 10226 -1296 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 -1296 10226
rect -1916 10102 -1296 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 -1296 10102
rect -1916 9978 -1296 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 -1296 9978
rect -1916 -1120 -1296 9922
rect -956 597212 -336 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 -336 597212
rect -956 597088 -336 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 -336 597088
rect -956 596964 -336 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 -336 596964
rect -956 596840 -336 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 -336 596840
rect -956 580350 -336 596784
rect 5418 597212 6038 598268
rect 5418 597156 5514 597212
rect 5570 597156 5638 597212
rect 5694 597156 5762 597212
rect 5818 597156 5886 597212
rect 5942 597156 6038 597212
rect 5418 597088 6038 597156
rect 5418 597032 5514 597088
rect 5570 597032 5638 597088
rect 5694 597032 5762 597088
rect 5818 597032 5886 597088
rect 5942 597032 6038 597088
rect 5418 596964 6038 597032
rect 5418 596908 5514 596964
rect 5570 596908 5638 596964
rect 5694 596908 5762 596964
rect 5818 596908 5886 596964
rect 5942 596908 6038 596964
rect 5418 596840 6038 596908
rect 5418 596784 5514 596840
rect 5570 596784 5638 596840
rect 5694 596784 5762 596840
rect 5818 596784 5886 596840
rect 5942 596784 6038 596840
rect -956 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 -336 580350
rect -956 580226 -336 580294
rect -956 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 -336 580226
rect -956 580102 -336 580170
rect -956 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 -336 580102
rect -956 579978 -336 580046
rect -956 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 -336 579978
rect -956 562350 -336 579922
rect 4172 587188 4228 587198
rect 4172 565124 4228 587132
rect 5418 580350 6038 596784
rect 9138 598172 9758 598268
rect 9138 598116 9234 598172
rect 9290 598116 9358 598172
rect 9414 598116 9482 598172
rect 9538 598116 9606 598172
rect 9662 598116 9758 598172
rect 9138 598048 9758 598116
rect 9138 597992 9234 598048
rect 9290 597992 9358 598048
rect 9414 597992 9482 598048
rect 9538 597992 9606 598048
rect 9662 597992 9758 598048
rect 9138 597924 9758 597992
rect 9138 597868 9234 597924
rect 9290 597868 9358 597924
rect 9414 597868 9482 597924
rect 9538 597868 9606 597924
rect 9662 597868 9758 597924
rect 9138 597800 9758 597868
rect 9138 597744 9234 597800
rect 9290 597744 9358 597800
rect 9414 597744 9482 597800
rect 9538 597744 9606 597800
rect 9662 597744 9758 597800
rect 9138 586350 9758 597744
rect 9138 586294 9234 586350
rect 9290 586294 9358 586350
rect 9414 586294 9482 586350
rect 9538 586294 9606 586350
rect 9662 586294 9758 586350
rect 9138 586226 9758 586294
rect 9138 586170 9234 586226
rect 9290 586170 9358 586226
rect 9414 586170 9482 586226
rect 9538 586170 9606 586226
rect 9662 586170 9758 586226
rect 9138 586102 9758 586170
rect 9138 586046 9234 586102
rect 9290 586046 9358 586102
rect 9414 586046 9482 586102
rect 9538 586046 9606 586102
rect 9662 586046 9758 586102
rect 9138 585978 9758 586046
rect 9138 585922 9234 585978
rect 9290 585922 9358 585978
rect 9414 585922 9482 585978
rect 9538 585922 9606 585978
rect 9662 585922 9758 585978
rect 9138 584990 9758 585922
rect 39858 598172 40478 598268
rect 39858 598116 39954 598172
rect 40010 598116 40078 598172
rect 40134 598116 40202 598172
rect 40258 598116 40326 598172
rect 40382 598116 40478 598172
rect 39858 598048 40478 598116
rect 39858 597992 39954 598048
rect 40010 597992 40078 598048
rect 40134 597992 40202 598048
rect 40258 597992 40326 598048
rect 40382 597992 40478 598048
rect 39858 597924 40478 597992
rect 39858 597868 39954 597924
rect 40010 597868 40078 597924
rect 40134 597868 40202 597924
rect 40258 597868 40326 597924
rect 40382 597868 40478 597924
rect 39858 597800 40478 597868
rect 39858 597744 39954 597800
rect 40010 597744 40078 597800
rect 40134 597744 40202 597800
rect 40258 597744 40326 597800
rect 40382 597744 40478 597800
rect 39858 586350 40478 597744
rect 39858 586294 39954 586350
rect 40010 586294 40078 586350
rect 40134 586294 40202 586350
rect 40258 586294 40326 586350
rect 40382 586294 40478 586350
rect 39858 586226 40478 586294
rect 39858 586170 39954 586226
rect 40010 586170 40078 586226
rect 40134 586170 40202 586226
rect 40258 586170 40326 586226
rect 40382 586170 40478 586226
rect 39858 586102 40478 586170
rect 39858 586046 39954 586102
rect 40010 586046 40078 586102
rect 40134 586046 40202 586102
rect 40258 586046 40326 586102
rect 40382 586046 40478 586102
rect 39858 585978 40478 586046
rect 39858 585922 39954 585978
rect 40010 585922 40078 585978
rect 40134 585922 40202 585978
rect 40258 585922 40326 585978
rect 40382 585922 40478 585978
rect 39858 584990 40478 585922
rect 70578 598172 71198 598268
rect 70578 598116 70674 598172
rect 70730 598116 70798 598172
rect 70854 598116 70922 598172
rect 70978 598116 71046 598172
rect 71102 598116 71198 598172
rect 70578 598048 71198 598116
rect 70578 597992 70674 598048
rect 70730 597992 70798 598048
rect 70854 597992 70922 598048
rect 70978 597992 71046 598048
rect 71102 597992 71198 598048
rect 70578 597924 71198 597992
rect 70578 597868 70674 597924
rect 70730 597868 70798 597924
rect 70854 597868 70922 597924
rect 70978 597868 71046 597924
rect 71102 597868 71198 597924
rect 70578 597800 71198 597868
rect 70578 597744 70674 597800
rect 70730 597744 70798 597800
rect 70854 597744 70922 597800
rect 70978 597744 71046 597800
rect 71102 597744 71198 597800
rect 70578 586350 71198 597744
rect 70578 586294 70674 586350
rect 70730 586294 70798 586350
rect 70854 586294 70922 586350
rect 70978 586294 71046 586350
rect 71102 586294 71198 586350
rect 70578 586226 71198 586294
rect 70578 586170 70674 586226
rect 70730 586170 70798 586226
rect 70854 586170 70922 586226
rect 70978 586170 71046 586226
rect 71102 586170 71198 586226
rect 70578 586102 71198 586170
rect 70578 586046 70674 586102
rect 70730 586046 70798 586102
rect 70854 586046 70922 586102
rect 70978 586046 71046 586102
rect 71102 586046 71198 586102
rect 70578 585978 71198 586046
rect 70578 585922 70674 585978
rect 70730 585922 70798 585978
rect 70854 585922 70922 585978
rect 70978 585922 71046 585978
rect 71102 585922 71198 585978
rect 70578 584990 71198 585922
rect 101298 598172 101918 598268
rect 101298 598116 101394 598172
rect 101450 598116 101518 598172
rect 101574 598116 101642 598172
rect 101698 598116 101766 598172
rect 101822 598116 101918 598172
rect 101298 598048 101918 598116
rect 101298 597992 101394 598048
rect 101450 597992 101518 598048
rect 101574 597992 101642 598048
rect 101698 597992 101766 598048
rect 101822 597992 101918 598048
rect 101298 597924 101918 597992
rect 101298 597868 101394 597924
rect 101450 597868 101518 597924
rect 101574 597868 101642 597924
rect 101698 597868 101766 597924
rect 101822 597868 101918 597924
rect 101298 597800 101918 597868
rect 101298 597744 101394 597800
rect 101450 597744 101518 597800
rect 101574 597744 101642 597800
rect 101698 597744 101766 597800
rect 101822 597744 101918 597800
rect 101298 586350 101918 597744
rect 101298 586294 101394 586350
rect 101450 586294 101518 586350
rect 101574 586294 101642 586350
rect 101698 586294 101766 586350
rect 101822 586294 101918 586350
rect 101298 586226 101918 586294
rect 101298 586170 101394 586226
rect 101450 586170 101518 586226
rect 101574 586170 101642 586226
rect 101698 586170 101766 586226
rect 101822 586170 101918 586226
rect 101298 586102 101918 586170
rect 101298 586046 101394 586102
rect 101450 586046 101518 586102
rect 101574 586046 101642 586102
rect 101698 586046 101766 586102
rect 101822 586046 101918 586102
rect 101298 585978 101918 586046
rect 101298 585922 101394 585978
rect 101450 585922 101518 585978
rect 101574 585922 101642 585978
rect 101698 585922 101766 585978
rect 101822 585922 101918 585978
rect 101298 584990 101918 585922
rect 132018 598172 132638 598268
rect 132018 598116 132114 598172
rect 132170 598116 132238 598172
rect 132294 598116 132362 598172
rect 132418 598116 132486 598172
rect 132542 598116 132638 598172
rect 132018 598048 132638 598116
rect 132018 597992 132114 598048
rect 132170 597992 132238 598048
rect 132294 597992 132362 598048
rect 132418 597992 132486 598048
rect 132542 597992 132638 598048
rect 132018 597924 132638 597992
rect 132018 597868 132114 597924
rect 132170 597868 132238 597924
rect 132294 597868 132362 597924
rect 132418 597868 132486 597924
rect 132542 597868 132638 597924
rect 132018 597800 132638 597868
rect 132018 597744 132114 597800
rect 132170 597744 132238 597800
rect 132294 597744 132362 597800
rect 132418 597744 132486 597800
rect 132542 597744 132638 597800
rect 132018 586350 132638 597744
rect 132018 586294 132114 586350
rect 132170 586294 132238 586350
rect 132294 586294 132362 586350
rect 132418 586294 132486 586350
rect 132542 586294 132638 586350
rect 132018 586226 132638 586294
rect 132018 586170 132114 586226
rect 132170 586170 132238 586226
rect 132294 586170 132362 586226
rect 132418 586170 132486 586226
rect 132542 586170 132638 586226
rect 132018 586102 132638 586170
rect 132018 586046 132114 586102
rect 132170 586046 132238 586102
rect 132294 586046 132362 586102
rect 132418 586046 132486 586102
rect 132542 586046 132638 586102
rect 132018 585978 132638 586046
rect 132018 585922 132114 585978
rect 132170 585922 132238 585978
rect 132294 585922 132362 585978
rect 132418 585922 132486 585978
rect 132542 585922 132638 585978
rect 132018 584990 132638 585922
rect 162738 598172 163358 598268
rect 162738 598116 162834 598172
rect 162890 598116 162958 598172
rect 163014 598116 163082 598172
rect 163138 598116 163206 598172
rect 163262 598116 163358 598172
rect 162738 598048 163358 598116
rect 162738 597992 162834 598048
rect 162890 597992 162958 598048
rect 163014 597992 163082 598048
rect 163138 597992 163206 598048
rect 163262 597992 163358 598048
rect 162738 597924 163358 597992
rect 162738 597868 162834 597924
rect 162890 597868 162958 597924
rect 163014 597868 163082 597924
rect 163138 597868 163206 597924
rect 163262 597868 163358 597924
rect 162738 597800 163358 597868
rect 162738 597744 162834 597800
rect 162890 597744 162958 597800
rect 163014 597744 163082 597800
rect 163138 597744 163206 597800
rect 163262 597744 163358 597800
rect 162738 586350 163358 597744
rect 162738 586294 162834 586350
rect 162890 586294 162958 586350
rect 163014 586294 163082 586350
rect 163138 586294 163206 586350
rect 163262 586294 163358 586350
rect 162738 586226 163358 586294
rect 162738 586170 162834 586226
rect 162890 586170 162958 586226
rect 163014 586170 163082 586226
rect 163138 586170 163206 586226
rect 163262 586170 163358 586226
rect 162738 586102 163358 586170
rect 162738 586046 162834 586102
rect 162890 586046 162958 586102
rect 163014 586046 163082 586102
rect 163138 586046 163206 586102
rect 163262 586046 163358 586102
rect 162738 585978 163358 586046
rect 162738 585922 162834 585978
rect 162890 585922 162958 585978
rect 163014 585922 163082 585978
rect 163138 585922 163206 585978
rect 163262 585922 163358 585978
rect 162738 584990 163358 585922
rect 193458 598172 194078 598268
rect 193458 598116 193554 598172
rect 193610 598116 193678 598172
rect 193734 598116 193802 598172
rect 193858 598116 193926 598172
rect 193982 598116 194078 598172
rect 193458 598048 194078 598116
rect 193458 597992 193554 598048
rect 193610 597992 193678 598048
rect 193734 597992 193802 598048
rect 193858 597992 193926 598048
rect 193982 597992 194078 598048
rect 193458 597924 194078 597992
rect 193458 597868 193554 597924
rect 193610 597868 193678 597924
rect 193734 597868 193802 597924
rect 193858 597868 193926 597924
rect 193982 597868 194078 597924
rect 193458 597800 194078 597868
rect 193458 597744 193554 597800
rect 193610 597744 193678 597800
rect 193734 597744 193802 597800
rect 193858 597744 193926 597800
rect 193982 597744 194078 597800
rect 193458 586350 194078 597744
rect 193458 586294 193554 586350
rect 193610 586294 193678 586350
rect 193734 586294 193802 586350
rect 193858 586294 193926 586350
rect 193982 586294 194078 586350
rect 193458 586226 194078 586294
rect 193458 586170 193554 586226
rect 193610 586170 193678 586226
rect 193734 586170 193802 586226
rect 193858 586170 193926 586226
rect 193982 586170 194078 586226
rect 193458 586102 194078 586170
rect 193458 586046 193554 586102
rect 193610 586046 193678 586102
rect 193734 586046 193802 586102
rect 193858 586046 193926 586102
rect 193982 586046 194078 586102
rect 193458 585978 194078 586046
rect 193458 585922 193554 585978
rect 193610 585922 193678 585978
rect 193734 585922 193802 585978
rect 193858 585922 193926 585978
rect 193982 585922 194078 585978
rect 193458 584990 194078 585922
rect 224178 598172 224798 598268
rect 224178 598116 224274 598172
rect 224330 598116 224398 598172
rect 224454 598116 224522 598172
rect 224578 598116 224646 598172
rect 224702 598116 224798 598172
rect 224178 598048 224798 598116
rect 224178 597992 224274 598048
rect 224330 597992 224398 598048
rect 224454 597992 224522 598048
rect 224578 597992 224646 598048
rect 224702 597992 224798 598048
rect 224178 597924 224798 597992
rect 224178 597868 224274 597924
rect 224330 597868 224398 597924
rect 224454 597868 224522 597924
rect 224578 597868 224646 597924
rect 224702 597868 224798 597924
rect 224178 597800 224798 597868
rect 224178 597744 224274 597800
rect 224330 597744 224398 597800
rect 224454 597744 224522 597800
rect 224578 597744 224646 597800
rect 224702 597744 224798 597800
rect 224178 586350 224798 597744
rect 224178 586294 224274 586350
rect 224330 586294 224398 586350
rect 224454 586294 224522 586350
rect 224578 586294 224646 586350
rect 224702 586294 224798 586350
rect 224178 586226 224798 586294
rect 224178 586170 224274 586226
rect 224330 586170 224398 586226
rect 224454 586170 224522 586226
rect 224578 586170 224646 586226
rect 224702 586170 224798 586226
rect 224178 586102 224798 586170
rect 224178 586046 224274 586102
rect 224330 586046 224398 586102
rect 224454 586046 224522 586102
rect 224578 586046 224646 586102
rect 224702 586046 224798 586102
rect 224178 585978 224798 586046
rect 224178 585922 224274 585978
rect 224330 585922 224398 585978
rect 224454 585922 224522 585978
rect 224578 585922 224646 585978
rect 224702 585922 224798 585978
rect 224178 584990 224798 585922
rect 254898 598172 255518 598268
rect 254898 598116 254994 598172
rect 255050 598116 255118 598172
rect 255174 598116 255242 598172
rect 255298 598116 255366 598172
rect 255422 598116 255518 598172
rect 254898 598048 255518 598116
rect 254898 597992 254994 598048
rect 255050 597992 255118 598048
rect 255174 597992 255242 598048
rect 255298 597992 255366 598048
rect 255422 597992 255518 598048
rect 254898 597924 255518 597992
rect 254898 597868 254994 597924
rect 255050 597868 255118 597924
rect 255174 597868 255242 597924
rect 255298 597868 255366 597924
rect 255422 597868 255518 597924
rect 254898 597800 255518 597868
rect 254898 597744 254994 597800
rect 255050 597744 255118 597800
rect 255174 597744 255242 597800
rect 255298 597744 255366 597800
rect 255422 597744 255518 597800
rect 254898 586350 255518 597744
rect 254898 586294 254994 586350
rect 255050 586294 255118 586350
rect 255174 586294 255242 586350
rect 255298 586294 255366 586350
rect 255422 586294 255518 586350
rect 254898 586226 255518 586294
rect 254898 586170 254994 586226
rect 255050 586170 255118 586226
rect 255174 586170 255242 586226
rect 255298 586170 255366 586226
rect 255422 586170 255518 586226
rect 254898 586102 255518 586170
rect 254898 586046 254994 586102
rect 255050 586046 255118 586102
rect 255174 586046 255242 586102
rect 255298 586046 255366 586102
rect 255422 586046 255518 586102
rect 254898 585978 255518 586046
rect 254898 585922 254994 585978
rect 255050 585922 255118 585978
rect 255174 585922 255242 585978
rect 255298 585922 255366 585978
rect 255422 585922 255518 585978
rect 254898 584990 255518 585922
rect 285618 598172 286238 598268
rect 285618 598116 285714 598172
rect 285770 598116 285838 598172
rect 285894 598116 285962 598172
rect 286018 598116 286086 598172
rect 286142 598116 286238 598172
rect 285618 598048 286238 598116
rect 285618 597992 285714 598048
rect 285770 597992 285838 598048
rect 285894 597992 285962 598048
rect 286018 597992 286086 598048
rect 286142 597992 286238 598048
rect 285618 597924 286238 597992
rect 285618 597868 285714 597924
rect 285770 597868 285838 597924
rect 285894 597868 285962 597924
rect 286018 597868 286086 597924
rect 286142 597868 286238 597924
rect 285618 597800 286238 597868
rect 285618 597744 285714 597800
rect 285770 597744 285838 597800
rect 285894 597744 285962 597800
rect 286018 597744 286086 597800
rect 286142 597744 286238 597800
rect 285618 586350 286238 597744
rect 285618 586294 285714 586350
rect 285770 586294 285838 586350
rect 285894 586294 285962 586350
rect 286018 586294 286086 586350
rect 286142 586294 286238 586350
rect 285618 586226 286238 586294
rect 285618 586170 285714 586226
rect 285770 586170 285838 586226
rect 285894 586170 285962 586226
rect 286018 586170 286086 586226
rect 286142 586170 286238 586226
rect 285618 586102 286238 586170
rect 285618 586046 285714 586102
rect 285770 586046 285838 586102
rect 285894 586046 285962 586102
rect 286018 586046 286086 586102
rect 286142 586046 286238 586102
rect 285618 585978 286238 586046
rect 285618 585922 285714 585978
rect 285770 585922 285838 585978
rect 285894 585922 285962 585978
rect 286018 585922 286086 585978
rect 286142 585922 286238 585978
rect 285618 584990 286238 585922
rect 316338 598172 316958 598268
rect 316338 598116 316434 598172
rect 316490 598116 316558 598172
rect 316614 598116 316682 598172
rect 316738 598116 316806 598172
rect 316862 598116 316958 598172
rect 316338 598048 316958 598116
rect 316338 597992 316434 598048
rect 316490 597992 316558 598048
rect 316614 597992 316682 598048
rect 316738 597992 316806 598048
rect 316862 597992 316958 598048
rect 316338 597924 316958 597992
rect 316338 597868 316434 597924
rect 316490 597868 316558 597924
rect 316614 597868 316682 597924
rect 316738 597868 316806 597924
rect 316862 597868 316958 597924
rect 316338 597800 316958 597868
rect 316338 597744 316434 597800
rect 316490 597744 316558 597800
rect 316614 597744 316682 597800
rect 316738 597744 316806 597800
rect 316862 597744 316958 597800
rect 316338 586350 316958 597744
rect 316338 586294 316434 586350
rect 316490 586294 316558 586350
rect 316614 586294 316682 586350
rect 316738 586294 316806 586350
rect 316862 586294 316958 586350
rect 316338 586226 316958 586294
rect 316338 586170 316434 586226
rect 316490 586170 316558 586226
rect 316614 586170 316682 586226
rect 316738 586170 316806 586226
rect 316862 586170 316958 586226
rect 316338 586102 316958 586170
rect 316338 586046 316434 586102
rect 316490 586046 316558 586102
rect 316614 586046 316682 586102
rect 316738 586046 316806 586102
rect 316862 586046 316958 586102
rect 316338 585978 316958 586046
rect 316338 585922 316434 585978
rect 316490 585922 316558 585978
rect 316614 585922 316682 585978
rect 316738 585922 316806 585978
rect 316862 585922 316958 585978
rect 316338 584990 316958 585922
rect 347058 598172 347678 598268
rect 347058 598116 347154 598172
rect 347210 598116 347278 598172
rect 347334 598116 347402 598172
rect 347458 598116 347526 598172
rect 347582 598116 347678 598172
rect 347058 598048 347678 598116
rect 347058 597992 347154 598048
rect 347210 597992 347278 598048
rect 347334 597992 347402 598048
rect 347458 597992 347526 598048
rect 347582 597992 347678 598048
rect 347058 597924 347678 597992
rect 347058 597868 347154 597924
rect 347210 597868 347278 597924
rect 347334 597868 347402 597924
rect 347458 597868 347526 597924
rect 347582 597868 347678 597924
rect 347058 597800 347678 597868
rect 347058 597744 347154 597800
rect 347210 597744 347278 597800
rect 347334 597744 347402 597800
rect 347458 597744 347526 597800
rect 347582 597744 347678 597800
rect 347058 586350 347678 597744
rect 347058 586294 347154 586350
rect 347210 586294 347278 586350
rect 347334 586294 347402 586350
rect 347458 586294 347526 586350
rect 347582 586294 347678 586350
rect 347058 586226 347678 586294
rect 347058 586170 347154 586226
rect 347210 586170 347278 586226
rect 347334 586170 347402 586226
rect 347458 586170 347526 586226
rect 347582 586170 347678 586226
rect 347058 586102 347678 586170
rect 347058 586046 347154 586102
rect 347210 586046 347278 586102
rect 347334 586046 347402 586102
rect 347458 586046 347526 586102
rect 347582 586046 347678 586102
rect 347058 585978 347678 586046
rect 347058 585922 347154 585978
rect 347210 585922 347278 585978
rect 347334 585922 347402 585978
rect 347458 585922 347526 585978
rect 347582 585922 347678 585978
rect 347058 584990 347678 585922
rect 377778 598172 378398 598268
rect 377778 598116 377874 598172
rect 377930 598116 377998 598172
rect 378054 598116 378122 598172
rect 378178 598116 378246 598172
rect 378302 598116 378398 598172
rect 377778 598048 378398 598116
rect 377778 597992 377874 598048
rect 377930 597992 377998 598048
rect 378054 597992 378122 598048
rect 378178 597992 378246 598048
rect 378302 597992 378398 598048
rect 377778 597924 378398 597992
rect 377778 597868 377874 597924
rect 377930 597868 377998 597924
rect 378054 597868 378122 597924
rect 378178 597868 378246 597924
rect 378302 597868 378398 597924
rect 377778 597800 378398 597868
rect 377778 597744 377874 597800
rect 377930 597744 377998 597800
rect 378054 597744 378122 597800
rect 378178 597744 378246 597800
rect 378302 597744 378398 597800
rect 377778 586350 378398 597744
rect 377778 586294 377874 586350
rect 377930 586294 377998 586350
rect 378054 586294 378122 586350
rect 378178 586294 378246 586350
rect 378302 586294 378398 586350
rect 377778 586226 378398 586294
rect 377778 586170 377874 586226
rect 377930 586170 377998 586226
rect 378054 586170 378122 586226
rect 378178 586170 378246 586226
rect 378302 586170 378398 586226
rect 377778 586102 378398 586170
rect 377778 586046 377874 586102
rect 377930 586046 377998 586102
rect 378054 586046 378122 586102
rect 378178 586046 378246 586102
rect 378302 586046 378398 586102
rect 377778 585978 378398 586046
rect 377778 585922 377874 585978
rect 377930 585922 377998 585978
rect 378054 585922 378122 585978
rect 378178 585922 378246 585978
rect 378302 585922 378398 585978
rect 377778 584990 378398 585922
rect 408498 598172 409118 598268
rect 408498 598116 408594 598172
rect 408650 598116 408718 598172
rect 408774 598116 408842 598172
rect 408898 598116 408966 598172
rect 409022 598116 409118 598172
rect 408498 598048 409118 598116
rect 408498 597992 408594 598048
rect 408650 597992 408718 598048
rect 408774 597992 408842 598048
rect 408898 597992 408966 598048
rect 409022 597992 409118 598048
rect 408498 597924 409118 597992
rect 408498 597868 408594 597924
rect 408650 597868 408718 597924
rect 408774 597868 408842 597924
rect 408898 597868 408966 597924
rect 409022 597868 409118 597924
rect 408498 597800 409118 597868
rect 408498 597744 408594 597800
rect 408650 597744 408718 597800
rect 408774 597744 408842 597800
rect 408898 597744 408966 597800
rect 409022 597744 409118 597800
rect 408498 586350 409118 597744
rect 408498 586294 408594 586350
rect 408650 586294 408718 586350
rect 408774 586294 408842 586350
rect 408898 586294 408966 586350
rect 409022 586294 409118 586350
rect 408498 586226 409118 586294
rect 408498 586170 408594 586226
rect 408650 586170 408718 586226
rect 408774 586170 408842 586226
rect 408898 586170 408966 586226
rect 409022 586170 409118 586226
rect 408498 586102 409118 586170
rect 408498 586046 408594 586102
rect 408650 586046 408718 586102
rect 408774 586046 408842 586102
rect 408898 586046 408966 586102
rect 409022 586046 409118 586102
rect 408498 585978 409118 586046
rect 408498 585922 408594 585978
rect 408650 585922 408718 585978
rect 408774 585922 408842 585978
rect 408898 585922 408966 585978
rect 409022 585922 409118 585978
rect 408498 584990 409118 585922
rect 439218 598172 439838 598268
rect 439218 598116 439314 598172
rect 439370 598116 439438 598172
rect 439494 598116 439562 598172
rect 439618 598116 439686 598172
rect 439742 598116 439838 598172
rect 439218 598048 439838 598116
rect 439218 597992 439314 598048
rect 439370 597992 439438 598048
rect 439494 597992 439562 598048
rect 439618 597992 439686 598048
rect 439742 597992 439838 598048
rect 439218 597924 439838 597992
rect 439218 597868 439314 597924
rect 439370 597868 439438 597924
rect 439494 597868 439562 597924
rect 439618 597868 439686 597924
rect 439742 597868 439838 597924
rect 439218 597800 439838 597868
rect 439218 597744 439314 597800
rect 439370 597744 439438 597800
rect 439494 597744 439562 597800
rect 439618 597744 439686 597800
rect 439742 597744 439838 597800
rect 439218 586350 439838 597744
rect 439218 586294 439314 586350
rect 439370 586294 439438 586350
rect 439494 586294 439562 586350
rect 439618 586294 439686 586350
rect 439742 586294 439838 586350
rect 439218 586226 439838 586294
rect 439218 586170 439314 586226
rect 439370 586170 439438 586226
rect 439494 586170 439562 586226
rect 439618 586170 439686 586226
rect 439742 586170 439838 586226
rect 439218 586102 439838 586170
rect 439218 586046 439314 586102
rect 439370 586046 439438 586102
rect 439494 586046 439562 586102
rect 439618 586046 439686 586102
rect 439742 586046 439838 586102
rect 439218 585978 439838 586046
rect 439218 585922 439314 585978
rect 439370 585922 439438 585978
rect 439494 585922 439562 585978
rect 439618 585922 439686 585978
rect 439742 585922 439838 585978
rect 439218 584990 439838 585922
rect 469938 598172 470558 598268
rect 469938 598116 470034 598172
rect 470090 598116 470158 598172
rect 470214 598116 470282 598172
rect 470338 598116 470406 598172
rect 470462 598116 470558 598172
rect 469938 598048 470558 598116
rect 469938 597992 470034 598048
rect 470090 597992 470158 598048
rect 470214 597992 470282 598048
rect 470338 597992 470406 598048
rect 470462 597992 470558 598048
rect 469938 597924 470558 597992
rect 469938 597868 470034 597924
rect 470090 597868 470158 597924
rect 470214 597868 470282 597924
rect 470338 597868 470406 597924
rect 470462 597868 470558 597924
rect 469938 597800 470558 597868
rect 469938 597744 470034 597800
rect 470090 597744 470158 597800
rect 470214 597744 470282 597800
rect 470338 597744 470406 597800
rect 470462 597744 470558 597800
rect 469938 586350 470558 597744
rect 469938 586294 470034 586350
rect 470090 586294 470158 586350
rect 470214 586294 470282 586350
rect 470338 586294 470406 586350
rect 470462 586294 470558 586350
rect 469938 586226 470558 586294
rect 469938 586170 470034 586226
rect 470090 586170 470158 586226
rect 470214 586170 470282 586226
rect 470338 586170 470406 586226
rect 470462 586170 470558 586226
rect 469938 586102 470558 586170
rect 469938 586046 470034 586102
rect 470090 586046 470158 586102
rect 470214 586046 470282 586102
rect 470338 586046 470406 586102
rect 470462 586046 470558 586102
rect 469938 585978 470558 586046
rect 469938 585922 470034 585978
rect 470090 585922 470158 585978
rect 470214 585922 470282 585978
rect 470338 585922 470406 585978
rect 470462 585922 470558 585978
rect 469938 584990 470558 585922
rect 500658 598172 501278 598268
rect 500658 598116 500754 598172
rect 500810 598116 500878 598172
rect 500934 598116 501002 598172
rect 501058 598116 501126 598172
rect 501182 598116 501278 598172
rect 500658 598048 501278 598116
rect 500658 597992 500754 598048
rect 500810 597992 500878 598048
rect 500934 597992 501002 598048
rect 501058 597992 501126 598048
rect 501182 597992 501278 598048
rect 500658 597924 501278 597992
rect 500658 597868 500754 597924
rect 500810 597868 500878 597924
rect 500934 597868 501002 597924
rect 501058 597868 501126 597924
rect 501182 597868 501278 597924
rect 500658 597800 501278 597868
rect 500658 597744 500754 597800
rect 500810 597744 500878 597800
rect 500934 597744 501002 597800
rect 501058 597744 501126 597800
rect 501182 597744 501278 597800
rect 500658 586350 501278 597744
rect 500658 586294 500754 586350
rect 500810 586294 500878 586350
rect 500934 586294 501002 586350
rect 501058 586294 501126 586350
rect 501182 586294 501278 586350
rect 500658 586226 501278 586294
rect 500658 586170 500754 586226
rect 500810 586170 500878 586226
rect 500934 586170 501002 586226
rect 501058 586170 501126 586226
rect 501182 586170 501278 586226
rect 500658 586102 501278 586170
rect 500658 586046 500754 586102
rect 500810 586046 500878 586102
rect 500934 586046 501002 586102
rect 501058 586046 501126 586102
rect 501182 586046 501278 586102
rect 500658 585978 501278 586046
rect 500658 585922 500754 585978
rect 500810 585922 500878 585978
rect 500934 585922 501002 585978
rect 501058 585922 501126 585978
rect 501182 585922 501278 585978
rect 500658 584990 501278 585922
rect 531378 598172 531998 598268
rect 531378 598116 531474 598172
rect 531530 598116 531598 598172
rect 531654 598116 531722 598172
rect 531778 598116 531846 598172
rect 531902 598116 531998 598172
rect 531378 598048 531998 598116
rect 531378 597992 531474 598048
rect 531530 597992 531598 598048
rect 531654 597992 531722 598048
rect 531778 597992 531846 598048
rect 531902 597992 531998 598048
rect 531378 597924 531998 597992
rect 531378 597868 531474 597924
rect 531530 597868 531598 597924
rect 531654 597868 531722 597924
rect 531778 597868 531846 597924
rect 531902 597868 531998 597924
rect 531378 597800 531998 597868
rect 531378 597744 531474 597800
rect 531530 597744 531598 597800
rect 531654 597744 531722 597800
rect 531778 597744 531846 597800
rect 531902 597744 531998 597800
rect 531378 586350 531998 597744
rect 531378 586294 531474 586350
rect 531530 586294 531598 586350
rect 531654 586294 531722 586350
rect 531778 586294 531846 586350
rect 531902 586294 531998 586350
rect 531378 586226 531998 586294
rect 531378 586170 531474 586226
rect 531530 586170 531598 586226
rect 531654 586170 531722 586226
rect 531778 586170 531846 586226
rect 531902 586170 531998 586226
rect 531378 586102 531998 586170
rect 531378 586046 531474 586102
rect 531530 586046 531598 586102
rect 531654 586046 531722 586102
rect 531778 586046 531846 586102
rect 531902 586046 531998 586102
rect 531378 585978 531998 586046
rect 531378 585922 531474 585978
rect 531530 585922 531598 585978
rect 531654 585922 531722 585978
rect 531778 585922 531846 585978
rect 531902 585922 531998 585978
rect 531378 584990 531998 585922
rect 562098 598172 562718 598268
rect 562098 598116 562194 598172
rect 562250 598116 562318 598172
rect 562374 598116 562442 598172
rect 562498 598116 562566 598172
rect 562622 598116 562718 598172
rect 562098 598048 562718 598116
rect 562098 597992 562194 598048
rect 562250 597992 562318 598048
rect 562374 597992 562442 598048
rect 562498 597992 562566 598048
rect 562622 597992 562718 598048
rect 562098 597924 562718 597992
rect 562098 597868 562194 597924
rect 562250 597868 562318 597924
rect 562374 597868 562442 597924
rect 562498 597868 562566 597924
rect 562622 597868 562718 597924
rect 562098 597800 562718 597868
rect 562098 597744 562194 597800
rect 562250 597744 562318 597800
rect 562374 597744 562442 597800
rect 562498 597744 562566 597800
rect 562622 597744 562718 597800
rect 562098 586350 562718 597744
rect 562098 586294 562194 586350
rect 562250 586294 562318 586350
rect 562374 586294 562442 586350
rect 562498 586294 562566 586350
rect 562622 586294 562718 586350
rect 562098 586226 562718 586294
rect 562098 586170 562194 586226
rect 562250 586170 562318 586226
rect 562374 586170 562442 586226
rect 562498 586170 562566 586226
rect 562622 586170 562718 586226
rect 562098 586102 562718 586170
rect 562098 586046 562194 586102
rect 562250 586046 562318 586102
rect 562374 586046 562442 586102
rect 562498 586046 562566 586102
rect 562622 586046 562718 586102
rect 562098 585978 562718 586046
rect 562098 585922 562194 585978
rect 562250 585922 562318 585978
rect 562374 585922 562442 585978
rect 562498 585922 562566 585978
rect 562622 585922 562718 585978
rect 562098 584990 562718 585922
rect 589098 597212 589718 598268
rect 589098 597156 589194 597212
rect 589250 597156 589318 597212
rect 589374 597156 589442 597212
rect 589498 597156 589566 597212
rect 589622 597156 589718 597212
rect 589098 597088 589718 597156
rect 589098 597032 589194 597088
rect 589250 597032 589318 597088
rect 589374 597032 589442 597088
rect 589498 597032 589566 597088
rect 589622 597032 589718 597088
rect 589098 596964 589718 597032
rect 589098 596908 589194 596964
rect 589250 596908 589318 596964
rect 589374 596908 589442 596964
rect 589498 596908 589566 596964
rect 589622 596908 589718 596964
rect 589098 596840 589718 596908
rect 589098 596784 589194 596840
rect 589250 596784 589318 596840
rect 589374 596784 589442 596840
rect 589498 596784 589566 596840
rect 589622 596784 589718 596840
rect 5418 580294 5514 580350
rect 5570 580294 5638 580350
rect 5694 580294 5762 580350
rect 5818 580294 5886 580350
rect 5942 580294 6038 580350
rect 5418 580226 6038 580294
rect 5418 580170 5514 580226
rect 5570 580170 5638 580226
rect 5694 580170 5762 580226
rect 5818 580170 5886 580226
rect 5942 580170 6038 580226
rect 5418 580102 6038 580170
rect 5418 580046 5514 580102
rect 5570 580046 5638 580102
rect 5694 580046 5762 580102
rect 5818 580046 5886 580102
rect 5942 580046 6038 580102
rect 5418 579978 6038 580046
rect 5418 579922 5514 579978
rect 5570 579922 5638 579978
rect 5694 579922 5762 579978
rect 5818 579922 5886 579978
rect 5942 579922 6038 579978
rect 4172 565058 4228 565068
rect 4284 573076 4340 573086
rect -956 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 -336 562350
rect -956 562226 -336 562294
rect -956 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 -336 562226
rect -956 562102 -336 562170
rect -956 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 -336 562102
rect -956 561978 -336 562046
rect -956 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 -336 561978
rect -956 544350 -336 561922
rect 4284 554596 4340 573020
rect 4284 554530 4340 554540
rect 5418 562350 6038 579922
rect 12448 580350 12768 580384
rect 12448 580294 12518 580350
rect 12574 580294 12642 580350
rect 12698 580294 12768 580350
rect 12448 580226 12768 580294
rect 12448 580170 12518 580226
rect 12574 580170 12642 580226
rect 12698 580170 12768 580226
rect 12448 580102 12768 580170
rect 12448 580046 12518 580102
rect 12574 580046 12642 580102
rect 12698 580046 12768 580102
rect 12448 579978 12768 580046
rect 12448 579922 12518 579978
rect 12574 579922 12642 579978
rect 12698 579922 12768 579978
rect 12448 579888 12768 579922
rect 43168 580350 43488 580384
rect 43168 580294 43238 580350
rect 43294 580294 43362 580350
rect 43418 580294 43488 580350
rect 43168 580226 43488 580294
rect 43168 580170 43238 580226
rect 43294 580170 43362 580226
rect 43418 580170 43488 580226
rect 43168 580102 43488 580170
rect 43168 580046 43238 580102
rect 43294 580046 43362 580102
rect 43418 580046 43488 580102
rect 43168 579978 43488 580046
rect 43168 579922 43238 579978
rect 43294 579922 43362 579978
rect 43418 579922 43488 579978
rect 43168 579888 43488 579922
rect 73888 580350 74208 580384
rect 73888 580294 73958 580350
rect 74014 580294 74082 580350
rect 74138 580294 74208 580350
rect 73888 580226 74208 580294
rect 73888 580170 73958 580226
rect 74014 580170 74082 580226
rect 74138 580170 74208 580226
rect 73888 580102 74208 580170
rect 73888 580046 73958 580102
rect 74014 580046 74082 580102
rect 74138 580046 74208 580102
rect 73888 579978 74208 580046
rect 73888 579922 73958 579978
rect 74014 579922 74082 579978
rect 74138 579922 74208 579978
rect 73888 579888 74208 579922
rect 104608 580350 104928 580384
rect 104608 580294 104678 580350
rect 104734 580294 104802 580350
rect 104858 580294 104928 580350
rect 104608 580226 104928 580294
rect 104608 580170 104678 580226
rect 104734 580170 104802 580226
rect 104858 580170 104928 580226
rect 104608 580102 104928 580170
rect 104608 580046 104678 580102
rect 104734 580046 104802 580102
rect 104858 580046 104928 580102
rect 104608 579978 104928 580046
rect 104608 579922 104678 579978
rect 104734 579922 104802 579978
rect 104858 579922 104928 579978
rect 104608 579888 104928 579922
rect 135328 580350 135648 580384
rect 135328 580294 135398 580350
rect 135454 580294 135522 580350
rect 135578 580294 135648 580350
rect 135328 580226 135648 580294
rect 135328 580170 135398 580226
rect 135454 580170 135522 580226
rect 135578 580170 135648 580226
rect 135328 580102 135648 580170
rect 135328 580046 135398 580102
rect 135454 580046 135522 580102
rect 135578 580046 135648 580102
rect 135328 579978 135648 580046
rect 135328 579922 135398 579978
rect 135454 579922 135522 579978
rect 135578 579922 135648 579978
rect 135328 579888 135648 579922
rect 166048 580350 166368 580384
rect 166048 580294 166118 580350
rect 166174 580294 166242 580350
rect 166298 580294 166368 580350
rect 166048 580226 166368 580294
rect 166048 580170 166118 580226
rect 166174 580170 166242 580226
rect 166298 580170 166368 580226
rect 166048 580102 166368 580170
rect 166048 580046 166118 580102
rect 166174 580046 166242 580102
rect 166298 580046 166368 580102
rect 166048 579978 166368 580046
rect 166048 579922 166118 579978
rect 166174 579922 166242 579978
rect 166298 579922 166368 579978
rect 166048 579888 166368 579922
rect 196768 580350 197088 580384
rect 196768 580294 196838 580350
rect 196894 580294 196962 580350
rect 197018 580294 197088 580350
rect 196768 580226 197088 580294
rect 196768 580170 196838 580226
rect 196894 580170 196962 580226
rect 197018 580170 197088 580226
rect 196768 580102 197088 580170
rect 196768 580046 196838 580102
rect 196894 580046 196962 580102
rect 197018 580046 197088 580102
rect 196768 579978 197088 580046
rect 196768 579922 196838 579978
rect 196894 579922 196962 579978
rect 197018 579922 197088 579978
rect 196768 579888 197088 579922
rect 227488 580350 227808 580384
rect 227488 580294 227558 580350
rect 227614 580294 227682 580350
rect 227738 580294 227808 580350
rect 227488 580226 227808 580294
rect 227488 580170 227558 580226
rect 227614 580170 227682 580226
rect 227738 580170 227808 580226
rect 227488 580102 227808 580170
rect 227488 580046 227558 580102
rect 227614 580046 227682 580102
rect 227738 580046 227808 580102
rect 227488 579978 227808 580046
rect 227488 579922 227558 579978
rect 227614 579922 227682 579978
rect 227738 579922 227808 579978
rect 227488 579888 227808 579922
rect 258208 580350 258528 580384
rect 258208 580294 258278 580350
rect 258334 580294 258402 580350
rect 258458 580294 258528 580350
rect 258208 580226 258528 580294
rect 258208 580170 258278 580226
rect 258334 580170 258402 580226
rect 258458 580170 258528 580226
rect 258208 580102 258528 580170
rect 258208 580046 258278 580102
rect 258334 580046 258402 580102
rect 258458 580046 258528 580102
rect 258208 579978 258528 580046
rect 258208 579922 258278 579978
rect 258334 579922 258402 579978
rect 258458 579922 258528 579978
rect 258208 579888 258528 579922
rect 288928 580350 289248 580384
rect 288928 580294 288998 580350
rect 289054 580294 289122 580350
rect 289178 580294 289248 580350
rect 288928 580226 289248 580294
rect 288928 580170 288998 580226
rect 289054 580170 289122 580226
rect 289178 580170 289248 580226
rect 288928 580102 289248 580170
rect 288928 580046 288998 580102
rect 289054 580046 289122 580102
rect 289178 580046 289248 580102
rect 288928 579978 289248 580046
rect 288928 579922 288998 579978
rect 289054 579922 289122 579978
rect 289178 579922 289248 579978
rect 288928 579888 289248 579922
rect 319648 580350 319968 580384
rect 319648 580294 319718 580350
rect 319774 580294 319842 580350
rect 319898 580294 319968 580350
rect 319648 580226 319968 580294
rect 319648 580170 319718 580226
rect 319774 580170 319842 580226
rect 319898 580170 319968 580226
rect 319648 580102 319968 580170
rect 319648 580046 319718 580102
rect 319774 580046 319842 580102
rect 319898 580046 319968 580102
rect 319648 579978 319968 580046
rect 319648 579922 319718 579978
rect 319774 579922 319842 579978
rect 319898 579922 319968 579978
rect 319648 579888 319968 579922
rect 350368 580350 350688 580384
rect 350368 580294 350438 580350
rect 350494 580294 350562 580350
rect 350618 580294 350688 580350
rect 350368 580226 350688 580294
rect 350368 580170 350438 580226
rect 350494 580170 350562 580226
rect 350618 580170 350688 580226
rect 350368 580102 350688 580170
rect 350368 580046 350438 580102
rect 350494 580046 350562 580102
rect 350618 580046 350688 580102
rect 350368 579978 350688 580046
rect 350368 579922 350438 579978
rect 350494 579922 350562 579978
rect 350618 579922 350688 579978
rect 350368 579888 350688 579922
rect 381088 580350 381408 580384
rect 381088 580294 381158 580350
rect 381214 580294 381282 580350
rect 381338 580294 381408 580350
rect 381088 580226 381408 580294
rect 381088 580170 381158 580226
rect 381214 580170 381282 580226
rect 381338 580170 381408 580226
rect 381088 580102 381408 580170
rect 381088 580046 381158 580102
rect 381214 580046 381282 580102
rect 381338 580046 381408 580102
rect 381088 579978 381408 580046
rect 381088 579922 381158 579978
rect 381214 579922 381282 579978
rect 381338 579922 381408 579978
rect 381088 579888 381408 579922
rect 411808 580350 412128 580384
rect 411808 580294 411878 580350
rect 411934 580294 412002 580350
rect 412058 580294 412128 580350
rect 411808 580226 412128 580294
rect 411808 580170 411878 580226
rect 411934 580170 412002 580226
rect 412058 580170 412128 580226
rect 411808 580102 412128 580170
rect 411808 580046 411878 580102
rect 411934 580046 412002 580102
rect 412058 580046 412128 580102
rect 411808 579978 412128 580046
rect 411808 579922 411878 579978
rect 411934 579922 412002 579978
rect 412058 579922 412128 579978
rect 411808 579888 412128 579922
rect 442528 580350 442848 580384
rect 442528 580294 442598 580350
rect 442654 580294 442722 580350
rect 442778 580294 442848 580350
rect 442528 580226 442848 580294
rect 442528 580170 442598 580226
rect 442654 580170 442722 580226
rect 442778 580170 442848 580226
rect 442528 580102 442848 580170
rect 442528 580046 442598 580102
rect 442654 580046 442722 580102
rect 442778 580046 442848 580102
rect 442528 579978 442848 580046
rect 442528 579922 442598 579978
rect 442654 579922 442722 579978
rect 442778 579922 442848 579978
rect 442528 579888 442848 579922
rect 473248 580350 473568 580384
rect 473248 580294 473318 580350
rect 473374 580294 473442 580350
rect 473498 580294 473568 580350
rect 473248 580226 473568 580294
rect 473248 580170 473318 580226
rect 473374 580170 473442 580226
rect 473498 580170 473568 580226
rect 473248 580102 473568 580170
rect 473248 580046 473318 580102
rect 473374 580046 473442 580102
rect 473498 580046 473568 580102
rect 473248 579978 473568 580046
rect 473248 579922 473318 579978
rect 473374 579922 473442 579978
rect 473498 579922 473568 579978
rect 473248 579888 473568 579922
rect 503968 580350 504288 580384
rect 503968 580294 504038 580350
rect 504094 580294 504162 580350
rect 504218 580294 504288 580350
rect 503968 580226 504288 580294
rect 503968 580170 504038 580226
rect 504094 580170 504162 580226
rect 504218 580170 504288 580226
rect 503968 580102 504288 580170
rect 503968 580046 504038 580102
rect 504094 580046 504162 580102
rect 504218 580046 504288 580102
rect 503968 579978 504288 580046
rect 503968 579922 504038 579978
rect 504094 579922 504162 579978
rect 504218 579922 504288 579978
rect 503968 579888 504288 579922
rect 534688 580350 535008 580384
rect 534688 580294 534758 580350
rect 534814 580294 534882 580350
rect 534938 580294 535008 580350
rect 534688 580226 535008 580294
rect 534688 580170 534758 580226
rect 534814 580170 534882 580226
rect 534938 580170 535008 580226
rect 534688 580102 535008 580170
rect 534688 580046 534758 580102
rect 534814 580046 534882 580102
rect 534938 580046 535008 580102
rect 534688 579978 535008 580046
rect 534688 579922 534758 579978
rect 534814 579922 534882 579978
rect 534938 579922 535008 579978
rect 534688 579888 535008 579922
rect 565408 580350 565728 580384
rect 565408 580294 565478 580350
rect 565534 580294 565602 580350
rect 565658 580294 565728 580350
rect 565408 580226 565728 580294
rect 565408 580170 565478 580226
rect 565534 580170 565602 580226
rect 565658 580170 565728 580226
rect 565408 580102 565728 580170
rect 565408 580046 565478 580102
rect 565534 580046 565602 580102
rect 565658 580046 565728 580102
rect 565408 579978 565728 580046
rect 565408 579922 565478 579978
rect 565534 579922 565602 579978
rect 565658 579922 565728 579978
rect 565408 579888 565728 579922
rect 589098 580350 589718 596784
rect 592818 598172 593438 598268
rect 592818 598116 592914 598172
rect 592970 598116 593038 598172
rect 593094 598116 593162 598172
rect 593218 598116 593286 598172
rect 593342 598116 593438 598172
rect 592818 598048 593438 598116
rect 592818 597992 592914 598048
rect 592970 597992 593038 598048
rect 593094 597992 593162 598048
rect 593218 597992 593286 598048
rect 593342 597992 593438 598048
rect 592818 597924 593438 597992
rect 592818 597868 592914 597924
rect 592970 597868 593038 597924
rect 593094 597868 593162 597924
rect 593218 597868 593286 597924
rect 593342 597868 593438 597924
rect 592818 597800 593438 597868
rect 592818 597744 592914 597800
rect 592970 597744 593038 597800
rect 593094 597744 593162 597800
rect 593218 597744 593286 597800
rect 593342 597744 593438 597800
rect 589098 580294 589194 580350
rect 589250 580294 589318 580350
rect 589374 580294 589442 580350
rect 589498 580294 589566 580350
rect 589622 580294 589718 580350
rect 589098 580226 589718 580294
rect 589098 580170 589194 580226
rect 589250 580170 589318 580226
rect 589374 580170 589442 580226
rect 589498 580170 589566 580226
rect 589622 580170 589718 580226
rect 589098 580102 589718 580170
rect 589098 580046 589194 580102
rect 589250 580046 589318 580102
rect 589374 580046 589442 580102
rect 589498 580046 589566 580102
rect 589622 580046 589718 580102
rect 589098 579978 589718 580046
rect 589098 579922 589194 579978
rect 589250 579922 589318 579978
rect 589374 579922 589442 579978
rect 589498 579922 589566 579978
rect 589622 579922 589718 579978
rect 27808 568350 28128 568384
rect 27808 568294 27878 568350
rect 27934 568294 28002 568350
rect 28058 568294 28128 568350
rect 27808 568226 28128 568294
rect 27808 568170 27878 568226
rect 27934 568170 28002 568226
rect 28058 568170 28128 568226
rect 27808 568102 28128 568170
rect 27808 568046 27878 568102
rect 27934 568046 28002 568102
rect 28058 568046 28128 568102
rect 27808 567978 28128 568046
rect 27808 567922 27878 567978
rect 27934 567922 28002 567978
rect 28058 567922 28128 567978
rect 27808 567888 28128 567922
rect 58528 568350 58848 568384
rect 58528 568294 58598 568350
rect 58654 568294 58722 568350
rect 58778 568294 58848 568350
rect 58528 568226 58848 568294
rect 58528 568170 58598 568226
rect 58654 568170 58722 568226
rect 58778 568170 58848 568226
rect 58528 568102 58848 568170
rect 58528 568046 58598 568102
rect 58654 568046 58722 568102
rect 58778 568046 58848 568102
rect 58528 567978 58848 568046
rect 58528 567922 58598 567978
rect 58654 567922 58722 567978
rect 58778 567922 58848 567978
rect 58528 567888 58848 567922
rect 89248 568350 89568 568384
rect 89248 568294 89318 568350
rect 89374 568294 89442 568350
rect 89498 568294 89568 568350
rect 89248 568226 89568 568294
rect 89248 568170 89318 568226
rect 89374 568170 89442 568226
rect 89498 568170 89568 568226
rect 89248 568102 89568 568170
rect 89248 568046 89318 568102
rect 89374 568046 89442 568102
rect 89498 568046 89568 568102
rect 89248 567978 89568 568046
rect 89248 567922 89318 567978
rect 89374 567922 89442 567978
rect 89498 567922 89568 567978
rect 89248 567888 89568 567922
rect 119968 568350 120288 568384
rect 119968 568294 120038 568350
rect 120094 568294 120162 568350
rect 120218 568294 120288 568350
rect 119968 568226 120288 568294
rect 119968 568170 120038 568226
rect 120094 568170 120162 568226
rect 120218 568170 120288 568226
rect 119968 568102 120288 568170
rect 119968 568046 120038 568102
rect 120094 568046 120162 568102
rect 120218 568046 120288 568102
rect 119968 567978 120288 568046
rect 119968 567922 120038 567978
rect 120094 567922 120162 567978
rect 120218 567922 120288 567978
rect 119968 567888 120288 567922
rect 150688 568350 151008 568384
rect 150688 568294 150758 568350
rect 150814 568294 150882 568350
rect 150938 568294 151008 568350
rect 150688 568226 151008 568294
rect 150688 568170 150758 568226
rect 150814 568170 150882 568226
rect 150938 568170 151008 568226
rect 150688 568102 151008 568170
rect 150688 568046 150758 568102
rect 150814 568046 150882 568102
rect 150938 568046 151008 568102
rect 150688 567978 151008 568046
rect 150688 567922 150758 567978
rect 150814 567922 150882 567978
rect 150938 567922 151008 567978
rect 150688 567888 151008 567922
rect 181408 568350 181728 568384
rect 181408 568294 181478 568350
rect 181534 568294 181602 568350
rect 181658 568294 181728 568350
rect 181408 568226 181728 568294
rect 181408 568170 181478 568226
rect 181534 568170 181602 568226
rect 181658 568170 181728 568226
rect 181408 568102 181728 568170
rect 181408 568046 181478 568102
rect 181534 568046 181602 568102
rect 181658 568046 181728 568102
rect 181408 567978 181728 568046
rect 181408 567922 181478 567978
rect 181534 567922 181602 567978
rect 181658 567922 181728 567978
rect 181408 567888 181728 567922
rect 212128 568350 212448 568384
rect 212128 568294 212198 568350
rect 212254 568294 212322 568350
rect 212378 568294 212448 568350
rect 212128 568226 212448 568294
rect 212128 568170 212198 568226
rect 212254 568170 212322 568226
rect 212378 568170 212448 568226
rect 212128 568102 212448 568170
rect 212128 568046 212198 568102
rect 212254 568046 212322 568102
rect 212378 568046 212448 568102
rect 212128 567978 212448 568046
rect 212128 567922 212198 567978
rect 212254 567922 212322 567978
rect 212378 567922 212448 567978
rect 212128 567888 212448 567922
rect 242848 568350 243168 568384
rect 242848 568294 242918 568350
rect 242974 568294 243042 568350
rect 243098 568294 243168 568350
rect 242848 568226 243168 568294
rect 242848 568170 242918 568226
rect 242974 568170 243042 568226
rect 243098 568170 243168 568226
rect 242848 568102 243168 568170
rect 242848 568046 242918 568102
rect 242974 568046 243042 568102
rect 243098 568046 243168 568102
rect 242848 567978 243168 568046
rect 242848 567922 242918 567978
rect 242974 567922 243042 567978
rect 243098 567922 243168 567978
rect 242848 567888 243168 567922
rect 273568 568350 273888 568384
rect 273568 568294 273638 568350
rect 273694 568294 273762 568350
rect 273818 568294 273888 568350
rect 273568 568226 273888 568294
rect 273568 568170 273638 568226
rect 273694 568170 273762 568226
rect 273818 568170 273888 568226
rect 273568 568102 273888 568170
rect 273568 568046 273638 568102
rect 273694 568046 273762 568102
rect 273818 568046 273888 568102
rect 273568 567978 273888 568046
rect 273568 567922 273638 567978
rect 273694 567922 273762 567978
rect 273818 567922 273888 567978
rect 273568 567888 273888 567922
rect 304288 568350 304608 568384
rect 304288 568294 304358 568350
rect 304414 568294 304482 568350
rect 304538 568294 304608 568350
rect 304288 568226 304608 568294
rect 304288 568170 304358 568226
rect 304414 568170 304482 568226
rect 304538 568170 304608 568226
rect 304288 568102 304608 568170
rect 304288 568046 304358 568102
rect 304414 568046 304482 568102
rect 304538 568046 304608 568102
rect 304288 567978 304608 568046
rect 304288 567922 304358 567978
rect 304414 567922 304482 567978
rect 304538 567922 304608 567978
rect 304288 567888 304608 567922
rect 335008 568350 335328 568384
rect 335008 568294 335078 568350
rect 335134 568294 335202 568350
rect 335258 568294 335328 568350
rect 335008 568226 335328 568294
rect 335008 568170 335078 568226
rect 335134 568170 335202 568226
rect 335258 568170 335328 568226
rect 335008 568102 335328 568170
rect 335008 568046 335078 568102
rect 335134 568046 335202 568102
rect 335258 568046 335328 568102
rect 335008 567978 335328 568046
rect 335008 567922 335078 567978
rect 335134 567922 335202 567978
rect 335258 567922 335328 567978
rect 335008 567888 335328 567922
rect 365728 568350 366048 568384
rect 365728 568294 365798 568350
rect 365854 568294 365922 568350
rect 365978 568294 366048 568350
rect 365728 568226 366048 568294
rect 365728 568170 365798 568226
rect 365854 568170 365922 568226
rect 365978 568170 366048 568226
rect 365728 568102 366048 568170
rect 365728 568046 365798 568102
rect 365854 568046 365922 568102
rect 365978 568046 366048 568102
rect 365728 567978 366048 568046
rect 365728 567922 365798 567978
rect 365854 567922 365922 567978
rect 365978 567922 366048 567978
rect 365728 567888 366048 567922
rect 396448 568350 396768 568384
rect 396448 568294 396518 568350
rect 396574 568294 396642 568350
rect 396698 568294 396768 568350
rect 396448 568226 396768 568294
rect 396448 568170 396518 568226
rect 396574 568170 396642 568226
rect 396698 568170 396768 568226
rect 396448 568102 396768 568170
rect 396448 568046 396518 568102
rect 396574 568046 396642 568102
rect 396698 568046 396768 568102
rect 396448 567978 396768 568046
rect 396448 567922 396518 567978
rect 396574 567922 396642 567978
rect 396698 567922 396768 567978
rect 396448 567888 396768 567922
rect 427168 568350 427488 568384
rect 427168 568294 427238 568350
rect 427294 568294 427362 568350
rect 427418 568294 427488 568350
rect 427168 568226 427488 568294
rect 427168 568170 427238 568226
rect 427294 568170 427362 568226
rect 427418 568170 427488 568226
rect 427168 568102 427488 568170
rect 427168 568046 427238 568102
rect 427294 568046 427362 568102
rect 427418 568046 427488 568102
rect 427168 567978 427488 568046
rect 427168 567922 427238 567978
rect 427294 567922 427362 567978
rect 427418 567922 427488 567978
rect 427168 567888 427488 567922
rect 457888 568350 458208 568384
rect 457888 568294 457958 568350
rect 458014 568294 458082 568350
rect 458138 568294 458208 568350
rect 457888 568226 458208 568294
rect 457888 568170 457958 568226
rect 458014 568170 458082 568226
rect 458138 568170 458208 568226
rect 457888 568102 458208 568170
rect 457888 568046 457958 568102
rect 458014 568046 458082 568102
rect 458138 568046 458208 568102
rect 457888 567978 458208 568046
rect 457888 567922 457958 567978
rect 458014 567922 458082 567978
rect 458138 567922 458208 567978
rect 457888 567888 458208 567922
rect 488608 568350 488928 568384
rect 488608 568294 488678 568350
rect 488734 568294 488802 568350
rect 488858 568294 488928 568350
rect 488608 568226 488928 568294
rect 488608 568170 488678 568226
rect 488734 568170 488802 568226
rect 488858 568170 488928 568226
rect 488608 568102 488928 568170
rect 488608 568046 488678 568102
rect 488734 568046 488802 568102
rect 488858 568046 488928 568102
rect 488608 567978 488928 568046
rect 488608 567922 488678 567978
rect 488734 567922 488802 567978
rect 488858 567922 488928 567978
rect 488608 567888 488928 567922
rect 519328 568350 519648 568384
rect 519328 568294 519398 568350
rect 519454 568294 519522 568350
rect 519578 568294 519648 568350
rect 519328 568226 519648 568294
rect 519328 568170 519398 568226
rect 519454 568170 519522 568226
rect 519578 568170 519648 568226
rect 519328 568102 519648 568170
rect 519328 568046 519398 568102
rect 519454 568046 519522 568102
rect 519578 568046 519648 568102
rect 519328 567978 519648 568046
rect 519328 567922 519398 567978
rect 519454 567922 519522 567978
rect 519578 567922 519648 567978
rect 519328 567888 519648 567922
rect 550048 568350 550368 568384
rect 550048 568294 550118 568350
rect 550174 568294 550242 568350
rect 550298 568294 550368 568350
rect 550048 568226 550368 568294
rect 550048 568170 550118 568226
rect 550174 568170 550242 568226
rect 550298 568170 550368 568226
rect 550048 568102 550368 568170
rect 550048 568046 550118 568102
rect 550174 568046 550242 568102
rect 550298 568046 550368 568102
rect 550048 567978 550368 568046
rect 550048 567922 550118 567978
rect 550174 567922 550242 567978
rect 550298 567922 550368 567978
rect 550048 567888 550368 567922
rect 5418 562294 5514 562350
rect 5570 562294 5638 562350
rect 5694 562294 5762 562350
rect 5818 562294 5886 562350
rect 5942 562294 6038 562350
rect 5418 562226 6038 562294
rect 5418 562170 5514 562226
rect 5570 562170 5638 562226
rect 5694 562170 5762 562226
rect 5818 562170 5886 562226
rect 5942 562170 6038 562226
rect 5418 562102 6038 562170
rect 5418 562046 5514 562102
rect 5570 562046 5638 562102
rect 5694 562046 5762 562102
rect 5818 562046 5886 562102
rect 5942 562046 6038 562102
rect 5418 561978 6038 562046
rect 5418 561922 5514 561978
rect 5570 561922 5638 561978
rect 5694 561922 5762 561978
rect 5818 561922 5886 561978
rect 5942 561922 6038 561978
rect -956 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 -336 544350
rect -956 544226 -336 544294
rect -956 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 -336 544226
rect -956 544102 -336 544170
rect -956 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 -336 544102
rect -956 543978 -336 544046
rect -956 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 -336 543978
rect -956 526350 -336 543922
rect -956 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 -336 526350
rect -956 526226 -336 526294
rect -956 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 -336 526226
rect -956 526102 -336 526170
rect -956 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 -336 526102
rect -956 525978 -336 526046
rect -956 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 -336 525978
rect -956 508350 -336 525922
rect 4172 544852 4228 544862
rect 4172 523012 4228 544796
rect 5418 544350 6038 561922
rect 12448 562350 12768 562384
rect 12448 562294 12518 562350
rect 12574 562294 12642 562350
rect 12698 562294 12768 562350
rect 12448 562226 12768 562294
rect 12448 562170 12518 562226
rect 12574 562170 12642 562226
rect 12698 562170 12768 562226
rect 12448 562102 12768 562170
rect 12448 562046 12518 562102
rect 12574 562046 12642 562102
rect 12698 562046 12768 562102
rect 12448 561978 12768 562046
rect 12448 561922 12518 561978
rect 12574 561922 12642 561978
rect 12698 561922 12768 561978
rect 12448 561888 12768 561922
rect 43168 562350 43488 562384
rect 43168 562294 43238 562350
rect 43294 562294 43362 562350
rect 43418 562294 43488 562350
rect 43168 562226 43488 562294
rect 43168 562170 43238 562226
rect 43294 562170 43362 562226
rect 43418 562170 43488 562226
rect 43168 562102 43488 562170
rect 43168 562046 43238 562102
rect 43294 562046 43362 562102
rect 43418 562046 43488 562102
rect 43168 561978 43488 562046
rect 43168 561922 43238 561978
rect 43294 561922 43362 561978
rect 43418 561922 43488 561978
rect 43168 561888 43488 561922
rect 73888 562350 74208 562384
rect 73888 562294 73958 562350
rect 74014 562294 74082 562350
rect 74138 562294 74208 562350
rect 73888 562226 74208 562294
rect 73888 562170 73958 562226
rect 74014 562170 74082 562226
rect 74138 562170 74208 562226
rect 73888 562102 74208 562170
rect 73888 562046 73958 562102
rect 74014 562046 74082 562102
rect 74138 562046 74208 562102
rect 73888 561978 74208 562046
rect 73888 561922 73958 561978
rect 74014 561922 74082 561978
rect 74138 561922 74208 561978
rect 73888 561888 74208 561922
rect 104608 562350 104928 562384
rect 104608 562294 104678 562350
rect 104734 562294 104802 562350
rect 104858 562294 104928 562350
rect 104608 562226 104928 562294
rect 104608 562170 104678 562226
rect 104734 562170 104802 562226
rect 104858 562170 104928 562226
rect 104608 562102 104928 562170
rect 104608 562046 104678 562102
rect 104734 562046 104802 562102
rect 104858 562046 104928 562102
rect 104608 561978 104928 562046
rect 104608 561922 104678 561978
rect 104734 561922 104802 561978
rect 104858 561922 104928 561978
rect 104608 561888 104928 561922
rect 135328 562350 135648 562384
rect 135328 562294 135398 562350
rect 135454 562294 135522 562350
rect 135578 562294 135648 562350
rect 135328 562226 135648 562294
rect 135328 562170 135398 562226
rect 135454 562170 135522 562226
rect 135578 562170 135648 562226
rect 135328 562102 135648 562170
rect 135328 562046 135398 562102
rect 135454 562046 135522 562102
rect 135578 562046 135648 562102
rect 135328 561978 135648 562046
rect 135328 561922 135398 561978
rect 135454 561922 135522 561978
rect 135578 561922 135648 561978
rect 135328 561888 135648 561922
rect 166048 562350 166368 562384
rect 166048 562294 166118 562350
rect 166174 562294 166242 562350
rect 166298 562294 166368 562350
rect 166048 562226 166368 562294
rect 166048 562170 166118 562226
rect 166174 562170 166242 562226
rect 166298 562170 166368 562226
rect 166048 562102 166368 562170
rect 166048 562046 166118 562102
rect 166174 562046 166242 562102
rect 166298 562046 166368 562102
rect 166048 561978 166368 562046
rect 166048 561922 166118 561978
rect 166174 561922 166242 561978
rect 166298 561922 166368 561978
rect 166048 561888 166368 561922
rect 196768 562350 197088 562384
rect 196768 562294 196838 562350
rect 196894 562294 196962 562350
rect 197018 562294 197088 562350
rect 196768 562226 197088 562294
rect 196768 562170 196838 562226
rect 196894 562170 196962 562226
rect 197018 562170 197088 562226
rect 196768 562102 197088 562170
rect 196768 562046 196838 562102
rect 196894 562046 196962 562102
rect 197018 562046 197088 562102
rect 196768 561978 197088 562046
rect 196768 561922 196838 561978
rect 196894 561922 196962 561978
rect 197018 561922 197088 561978
rect 196768 561888 197088 561922
rect 227488 562350 227808 562384
rect 227488 562294 227558 562350
rect 227614 562294 227682 562350
rect 227738 562294 227808 562350
rect 227488 562226 227808 562294
rect 227488 562170 227558 562226
rect 227614 562170 227682 562226
rect 227738 562170 227808 562226
rect 227488 562102 227808 562170
rect 227488 562046 227558 562102
rect 227614 562046 227682 562102
rect 227738 562046 227808 562102
rect 227488 561978 227808 562046
rect 227488 561922 227558 561978
rect 227614 561922 227682 561978
rect 227738 561922 227808 561978
rect 227488 561888 227808 561922
rect 258208 562350 258528 562384
rect 258208 562294 258278 562350
rect 258334 562294 258402 562350
rect 258458 562294 258528 562350
rect 258208 562226 258528 562294
rect 258208 562170 258278 562226
rect 258334 562170 258402 562226
rect 258458 562170 258528 562226
rect 258208 562102 258528 562170
rect 258208 562046 258278 562102
rect 258334 562046 258402 562102
rect 258458 562046 258528 562102
rect 258208 561978 258528 562046
rect 258208 561922 258278 561978
rect 258334 561922 258402 561978
rect 258458 561922 258528 561978
rect 258208 561888 258528 561922
rect 288928 562350 289248 562384
rect 288928 562294 288998 562350
rect 289054 562294 289122 562350
rect 289178 562294 289248 562350
rect 288928 562226 289248 562294
rect 288928 562170 288998 562226
rect 289054 562170 289122 562226
rect 289178 562170 289248 562226
rect 288928 562102 289248 562170
rect 288928 562046 288998 562102
rect 289054 562046 289122 562102
rect 289178 562046 289248 562102
rect 288928 561978 289248 562046
rect 288928 561922 288998 561978
rect 289054 561922 289122 561978
rect 289178 561922 289248 561978
rect 288928 561888 289248 561922
rect 319648 562350 319968 562384
rect 319648 562294 319718 562350
rect 319774 562294 319842 562350
rect 319898 562294 319968 562350
rect 319648 562226 319968 562294
rect 319648 562170 319718 562226
rect 319774 562170 319842 562226
rect 319898 562170 319968 562226
rect 319648 562102 319968 562170
rect 319648 562046 319718 562102
rect 319774 562046 319842 562102
rect 319898 562046 319968 562102
rect 319648 561978 319968 562046
rect 319648 561922 319718 561978
rect 319774 561922 319842 561978
rect 319898 561922 319968 561978
rect 319648 561888 319968 561922
rect 350368 562350 350688 562384
rect 350368 562294 350438 562350
rect 350494 562294 350562 562350
rect 350618 562294 350688 562350
rect 350368 562226 350688 562294
rect 350368 562170 350438 562226
rect 350494 562170 350562 562226
rect 350618 562170 350688 562226
rect 350368 562102 350688 562170
rect 350368 562046 350438 562102
rect 350494 562046 350562 562102
rect 350618 562046 350688 562102
rect 350368 561978 350688 562046
rect 350368 561922 350438 561978
rect 350494 561922 350562 561978
rect 350618 561922 350688 561978
rect 350368 561888 350688 561922
rect 381088 562350 381408 562384
rect 381088 562294 381158 562350
rect 381214 562294 381282 562350
rect 381338 562294 381408 562350
rect 381088 562226 381408 562294
rect 381088 562170 381158 562226
rect 381214 562170 381282 562226
rect 381338 562170 381408 562226
rect 381088 562102 381408 562170
rect 381088 562046 381158 562102
rect 381214 562046 381282 562102
rect 381338 562046 381408 562102
rect 381088 561978 381408 562046
rect 381088 561922 381158 561978
rect 381214 561922 381282 561978
rect 381338 561922 381408 561978
rect 381088 561888 381408 561922
rect 411808 562350 412128 562384
rect 411808 562294 411878 562350
rect 411934 562294 412002 562350
rect 412058 562294 412128 562350
rect 411808 562226 412128 562294
rect 411808 562170 411878 562226
rect 411934 562170 412002 562226
rect 412058 562170 412128 562226
rect 411808 562102 412128 562170
rect 411808 562046 411878 562102
rect 411934 562046 412002 562102
rect 412058 562046 412128 562102
rect 411808 561978 412128 562046
rect 411808 561922 411878 561978
rect 411934 561922 412002 561978
rect 412058 561922 412128 561978
rect 411808 561888 412128 561922
rect 442528 562350 442848 562384
rect 442528 562294 442598 562350
rect 442654 562294 442722 562350
rect 442778 562294 442848 562350
rect 442528 562226 442848 562294
rect 442528 562170 442598 562226
rect 442654 562170 442722 562226
rect 442778 562170 442848 562226
rect 442528 562102 442848 562170
rect 442528 562046 442598 562102
rect 442654 562046 442722 562102
rect 442778 562046 442848 562102
rect 442528 561978 442848 562046
rect 442528 561922 442598 561978
rect 442654 561922 442722 561978
rect 442778 561922 442848 561978
rect 442528 561888 442848 561922
rect 473248 562350 473568 562384
rect 473248 562294 473318 562350
rect 473374 562294 473442 562350
rect 473498 562294 473568 562350
rect 473248 562226 473568 562294
rect 473248 562170 473318 562226
rect 473374 562170 473442 562226
rect 473498 562170 473568 562226
rect 473248 562102 473568 562170
rect 473248 562046 473318 562102
rect 473374 562046 473442 562102
rect 473498 562046 473568 562102
rect 473248 561978 473568 562046
rect 473248 561922 473318 561978
rect 473374 561922 473442 561978
rect 473498 561922 473568 561978
rect 473248 561888 473568 561922
rect 503968 562350 504288 562384
rect 503968 562294 504038 562350
rect 504094 562294 504162 562350
rect 504218 562294 504288 562350
rect 503968 562226 504288 562294
rect 503968 562170 504038 562226
rect 504094 562170 504162 562226
rect 504218 562170 504288 562226
rect 503968 562102 504288 562170
rect 503968 562046 504038 562102
rect 504094 562046 504162 562102
rect 504218 562046 504288 562102
rect 503968 561978 504288 562046
rect 503968 561922 504038 561978
rect 504094 561922 504162 561978
rect 504218 561922 504288 561978
rect 503968 561888 504288 561922
rect 534688 562350 535008 562384
rect 534688 562294 534758 562350
rect 534814 562294 534882 562350
rect 534938 562294 535008 562350
rect 534688 562226 535008 562294
rect 534688 562170 534758 562226
rect 534814 562170 534882 562226
rect 534938 562170 535008 562226
rect 534688 562102 535008 562170
rect 534688 562046 534758 562102
rect 534814 562046 534882 562102
rect 534938 562046 535008 562102
rect 534688 561978 535008 562046
rect 534688 561922 534758 561978
rect 534814 561922 534882 561978
rect 534938 561922 535008 561978
rect 534688 561888 535008 561922
rect 565408 562350 565728 562384
rect 565408 562294 565478 562350
rect 565534 562294 565602 562350
rect 565658 562294 565728 562350
rect 565408 562226 565728 562294
rect 565408 562170 565478 562226
rect 565534 562170 565602 562226
rect 565658 562170 565728 562226
rect 589098 562350 589718 579922
rect 590492 588644 590548 588654
rect 590492 576324 590548 588588
rect 590492 576258 590548 576268
rect 592818 586350 593438 597744
rect 597360 598172 597980 598268
rect 597360 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect 597360 598048 597980 598116
rect 597360 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect 597360 597924 597980 597992
rect 597360 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect 597360 597800 597980 597868
rect 597360 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect 592818 586294 592914 586350
rect 592970 586294 593038 586350
rect 593094 586294 593162 586350
rect 593218 586294 593286 586350
rect 593342 586294 593438 586350
rect 592818 586226 593438 586294
rect 592818 586170 592914 586226
rect 592970 586170 593038 586226
rect 593094 586170 593162 586226
rect 593218 586170 593286 586226
rect 593342 586170 593438 586226
rect 592818 586102 593438 586170
rect 592818 586046 592914 586102
rect 592970 586046 593038 586102
rect 593094 586046 593162 586102
rect 593218 586046 593286 586102
rect 593342 586046 593438 586102
rect 592818 585978 593438 586046
rect 592818 585922 592914 585978
rect 592970 585922 593038 585978
rect 593094 585922 593162 585978
rect 593218 585922 593286 585978
rect 593342 585922 593438 585978
rect 591276 575428 591332 575438
rect 591276 565572 591332 575372
rect 591276 565506 591332 565516
rect 592818 568350 593438 585922
rect 592818 568294 592914 568350
rect 592970 568294 593038 568350
rect 593094 568294 593162 568350
rect 593218 568294 593286 568350
rect 593342 568294 593438 568350
rect 592818 568226 593438 568294
rect 592818 568170 592914 568226
rect 592970 568170 593038 568226
rect 593094 568170 593162 568226
rect 593218 568170 593286 568226
rect 593342 568170 593438 568226
rect 592818 568102 593438 568170
rect 592818 568046 592914 568102
rect 592970 568046 593038 568102
rect 593094 568046 593162 568102
rect 593218 568046 593286 568102
rect 593342 568046 593438 568102
rect 592818 567978 593438 568046
rect 592818 567922 592914 567978
rect 592970 567922 593038 567978
rect 593094 567922 593162 567978
rect 593218 567922 593286 567978
rect 593342 567922 593438 567978
rect 589098 562294 589194 562350
rect 589250 562294 589318 562350
rect 589374 562294 589442 562350
rect 589498 562294 589566 562350
rect 589622 562294 589718 562350
rect 589098 562226 589718 562294
rect 565408 562102 565728 562170
rect 565408 562046 565478 562102
rect 565534 562046 565602 562102
rect 565658 562046 565728 562102
rect 565408 561978 565728 562046
rect 565408 561922 565478 561978
rect 565534 561922 565602 561978
rect 565658 561922 565728 561978
rect 565408 561888 565728 561922
rect 586348 562212 586404 562222
rect 5418 544294 5514 544350
rect 5570 544294 5638 544350
rect 5694 544294 5762 544350
rect 5818 544294 5886 544350
rect 5942 544294 6038 544350
rect 5418 544226 6038 544294
rect 5418 544170 5514 544226
rect 5570 544170 5638 544226
rect 5694 544170 5762 544226
rect 5818 544170 5886 544226
rect 5942 544170 6038 544226
rect 5418 544102 6038 544170
rect 5418 544046 5514 544102
rect 5570 544046 5638 544102
rect 5694 544046 5762 544102
rect 5818 544046 5886 544102
rect 5942 544046 6038 544102
rect 5418 543978 6038 544046
rect 6188 558964 6244 558974
rect 6188 544068 6244 558908
rect 586348 554820 586404 562156
rect 586348 554754 586404 554764
rect 589098 562170 589194 562226
rect 589250 562170 589318 562226
rect 589374 562170 589442 562226
rect 589498 562170 589566 562226
rect 589622 562170 589718 562226
rect 589098 562102 589718 562170
rect 589098 562046 589194 562102
rect 589250 562046 589318 562102
rect 589374 562046 589442 562102
rect 589498 562046 589566 562102
rect 589622 562046 589718 562102
rect 589098 561978 589718 562046
rect 589098 561922 589194 561978
rect 589250 561922 589318 561978
rect 589374 561922 589442 561978
rect 589498 561922 589566 561978
rect 589622 561922 589718 561978
rect 27808 550350 28128 550384
rect 27808 550294 27878 550350
rect 27934 550294 28002 550350
rect 28058 550294 28128 550350
rect 27808 550226 28128 550294
rect 27808 550170 27878 550226
rect 27934 550170 28002 550226
rect 28058 550170 28128 550226
rect 27808 550102 28128 550170
rect 27808 550046 27878 550102
rect 27934 550046 28002 550102
rect 28058 550046 28128 550102
rect 27808 549978 28128 550046
rect 27808 549922 27878 549978
rect 27934 549922 28002 549978
rect 28058 549922 28128 549978
rect 27808 549888 28128 549922
rect 58528 550350 58848 550384
rect 58528 550294 58598 550350
rect 58654 550294 58722 550350
rect 58778 550294 58848 550350
rect 58528 550226 58848 550294
rect 58528 550170 58598 550226
rect 58654 550170 58722 550226
rect 58778 550170 58848 550226
rect 58528 550102 58848 550170
rect 58528 550046 58598 550102
rect 58654 550046 58722 550102
rect 58778 550046 58848 550102
rect 58528 549978 58848 550046
rect 58528 549922 58598 549978
rect 58654 549922 58722 549978
rect 58778 549922 58848 549978
rect 58528 549888 58848 549922
rect 89248 550350 89568 550384
rect 89248 550294 89318 550350
rect 89374 550294 89442 550350
rect 89498 550294 89568 550350
rect 89248 550226 89568 550294
rect 89248 550170 89318 550226
rect 89374 550170 89442 550226
rect 89498 550170 89568 550226
rect 89248 550102 89568 550170
rect 89248 550046 89318 550102
rect 89374 550046 89442 550102
rect 89498 550046 89568 550102
rect 89248 549978 89568 550046
rect 89248 549922 89318 549978
rect 89374 549922 89442 549978
rect 89498 549922 89568 549978
rect 89248 549888 89568 549922
rect 119968 550350 120288 550384
rect 119968 550294 120038 550350
rect 120094 550294 120162 550350
rect 120218 550294 120288 550350
rect 119968 550226 120288 550294
rect 119968 550170 120038 550226
rect 120094 550170 120162 550226
rect 120218 550170 120288 550226
rect 119968 550102 120288 550170
rect 119968 550046 120038 550102
rect 120094 550046 120162 550102
rect 120218 550046 120288 550102
rect 119968 549978 120288 550046
rect 119968 549922 120038 549978
rect 120094 549922 120162 549978
rect 120218 549922 120288 549978
rect 119968 549888 120288 549922
rect 150688 550350 151008 550384
rect 150688 550294 150758 550350
rect 150814 550294 150882 550350
rect 150938 550294 151008 550350
rect 150688 550226 151008 550294
rect 150688 550170 150758 550226
rect 150814 550170 150882 550226
rect 150938 550170 151008 550226
rect 150688 550102 151008 550170
rect 150688 550046 150758 550102
rect 150814 550046 150882 550102
rect 150938 550046 151008 550102
rect 150688 549978 151008 550046
rect 150688 549922 150758 549978
rect 150814 549922 150882 549978
rect 150938 549922 151008 549978
rect 150688 549888 151008 549922
rect 181408 550350 181728 550384
rect 181408 550294 181478 550350
rect 181534 550294 181602 550350
rect 181658 550294 181728 550350
rect 181408 550226 181728 550294
rect 181408 550170 181478 550226
rect 181534 550170 181602 550226
rect 181658 550170 181728 550226
rect 181408 550102 181728 550170
rect 181408 550046 181478 550102
rect 181534 550046 181602 550102
rect 181658 550046 181728 550102
rect 181408 549978 181728 550046
rect 181408 549922 181478 549978
rect 181534 549922 181602 549978
rect 181658 549922 181728 549978
rect 181408 549888 181728 549922
rect 212128 550350 212448 550384
rect 212128 550294 212198 550350
rect 212254 550294 212322 550350
rect 212378 550294 212448 550350
rect 212128 550226 212448 550294
rect 212128 550170 212198 550226
rect 212254 550170 212322 550226
rect 212378 550170 212448 550226
rect 212128 550102 212448 550170
rect 212128 550046 212198 550102
rect 212254 550046 212322 550102
rect 212378 550046 212448 550102
rect 212128 549978 212448 550046
rect 212128 549922 212198 549978
rect 212254 549922 212322 549978
rect 212378 549922 212448 549978
rect 212128 549888 212448 549922
rect 242848 550350 243168 550384
rect 242848 550294 242918 550350
rect 242974 550294 243042 550350
rect 243098 550294 243168 550350
rect 242848 550226 243168 550294
rect 242848 550170 242918 550226
rect 242974 550170 243042 550226
rect 243098 550170 243168 550226
rect 242848 550102 243168 550170
rect 242848 550046 242918 550102
rect 242974 550046 243042 550102
rect 243098 550046 243168 550102
rect 242848 549978 243168 550046
rect 242848 549922 242918 549978
rect 242974 549922 243042 549978
rect 243098 549922 243168 549978
rect 242848 549888 243168 549922
rect 273568 550350 273888 550384
rect 273568 550294 273638 550350
rect 273694 550294 273762 550350
rect 273818 550294 273888 550350
rect 273568 550226 273888 550294
rect 273568 550170 273638 550226
rect 273694 550170 273762 550226
rect 273818 550170 273888 550226
rect 273568 550102 273888 550170
rect 273568 550046 273638 550102
rect 273694 550046 273762 550102
rect 273818 550046 273888 550102
rect 273568 549978 273888 550046
rect 273568 549922 273638 549978
rect 273694 549922 273762 549978
rect 273818 549922 273888 549978
rect 273568 549888 273888 549922
rect 304288 550350 304608 550384
rect 304288 550294 304358 550350
rect 304414 550294 304482 550350
rect 304538 550294 304608 550350
rect 304288 550226 304608 550294
rect 304288 550170 304358 550226
rect 304414 550170 304482 550226
rect 304538 550170 304608 550226
rect 304288 550102 304608 550170
rect 304288 550046 304358 550102
rect 304414 550046 304482 550102
rect 304538 550046 304608 550102
rect 304288 549978 304608 550046
rect 304288 549922 304358 549978
rect 304414 549922 304482 549978
rect 304538 549922 304608 549978
rect 304288 549888 304608 549922
rect 335008 550350 335328 550384
rect 335008 550294 335078 550350
rect 335134 550294 335202 550350
rect 335258 550294 335328 550350
rect 335008 550226 335328 550294
rect 335008 550170 335078 550226
rect 335134 550170 335202 550226
rect 335258 550170 335328 550226
rect 335008 550102 335328 550170
rect 335008 550046 335078 550102
rect 335134 550046 335202 550102
rect 335258 550046 335328 550102
rect 335008 549978 335328 550046
rect 335008 549922 335078 549978
rect 335134 549922 335202 549978
rect 335258 549922 335328 549978
rect 335008 549888 335328 549922
rect 365728 550350 366048 550384
rect 365728 550294 365798 550350
rect 365854 550294 365922 550350
rect 365978 550294 366048 550350
rect 365728 550226 366048 550294
rect 365728 550170 365798 550226
rect 365854 550170 365922 550226
rect 365978 550170 366048 550226
rect 365728 550102 366048 550170
rect 365728 550046 365798 550102
rect 365854 550046 365922 550102
rect 365978 550046 366048 550102
rect 365728 549978 366048 550046
rect 365728 549922 365798 549978
rect 365854 549922 365922 549978
rect 365978 549922 366048 549978
rect 365728 549888 366048 549922
rect 396448 550350 396768 550384
rect 396448 550294 396518 550350
rect 396574 550294 396642 550350
rect 396698 550294 396768 550350
rect 396448 550226 396768 550294
rect 396448 550170 396518 550226
rect 396574 550170 396642 550226
rect 396698 550170 396768 550226
rect 396448 550102 396768 550170
rect 396448 550046 396518 550102
rect 396574 550046 396642 550102
rect 396698 550046 396768 550102
rect 396448 549978 396768 550046
rect 396448 549922 396518 549978
rect 396574 549922 396642 549978
rect 396698 549922 396768 549978
rect 396448 549888 396768 549922
rect 427168 550350 427488 550384
rect 427168 550294 427238 550350
rect 427294 550294 427362 550350
rect 427418 550294 427488 550350
rect 427168 550226 427488 550294
rect 427168 550170 427238 550226
rect 427294 550170 427362 550226
rect 427418 550170 427488 550226
rect 427168 550102 427488 550170
rect 427168 550046 427238 550102
rect 427294 550046 427362 550102
rect 427418 550046 427488 550102
rect 427168 549978 427488 550046
rect 427168 549922 427238 549978
rect 427294 549922 427362 549978
rect 427418 549922 427488 549978
rect 427168 549888 427488 549922
rect 457888 550350 458208 550384
rect 457888 550294 457958 550350
rect 458014 550294 458082 550350
rect 458138 550294 458208 550350
rect 457888 550226 458208 550294
rect 457888 550170 457958 550226
rect 458014 550170 458082 550226
rect 458138 550170 458208 550226
rect 457888 550102 458208 550170
rect 457888 550046 457958 550102
rect 458014 550046 458082 550102
rect 458138 550046 458208 550102
rect 457888 549978 458208 550046
rect 457888 549922 457958 549978
rect 458014 549922 458082 549978
rect 458138 549922 458208 549978
rect 457888 549888 458208 549922
rect 488608 550350 488928 550384
rect 488608 550294 488678 550350
rect 488734 550294 488802 550350
rect 488858 550294 488928 550350
rect 488608 550226 488928 550294
rect 488608 550170 488678 550226
rect 488734 550170 488802 550226
rect 488858 550170 488928 550226
rect 488608 550102 488928 550170
rect 488608 550046 488678 550102
rect 488734 550046 488802 550102
rect 488858 550046 488928 550102
rect 488608 549978 488928 550046
rect 488608 549922 488678 549978
rect 488734 549922 488802 549978
rect 488858 549922 488928 549978
rect 488608 549888 488928 549922
rect 519328 550350 519648 550384
rect 519328 550294 519398 550350
rect 519454 550294 519522 550350
rect 519578 550294 519648 550350
rect 519328 550226 519648 550294
rect 519328 550170 519398 550226
rect 519454 550170 519522 550226
rect 519578 550170 519648 550226
rect 519328 550102 519648 550170
rect 519328 550046 519398 550102
rect 519454 550046 519522 550102
rect 519578 550046 519648 550102
rect 519328 549978 519648 550046
rect 519328 549922 519398 549978
rect 519454 549922 519522 549978
rect 519578 549922 519648 549978
rect 519328 549888 519648 549922
rect 550048 550350 550368 550384
rect 550048 550294 550118 550350
rect 550174 550294 550242 550350
rect 550298 550294 550368 550350
rect 550048 550226 550368 550294
rect 550048 550170 550118 550226
rect 550174 550170 550242 550226
rect 550298 550170 550368 550226
rect 550048 550102 550368 550170
rect 550048 550046 550118 550102
rect 550174 550046 550242 550102
rect 550298 550046 550368 550102
rect 550048 549978 550368 550046
rect 550048 549922 550118 549978
rect 550174 549922 550242 549978
rect 550298 549922 550368 549978
rect 550048 549888 550368 549922
rect 6188 544002 6244 544012
rect 12448 544350 12768 544384
rect 12448 544294 12518 544350
rect 12574 544294 12642 544350
rect 12698 544294 12768 544350
rect 12448 544226 12768 544294
rect 12448 544170 12518 544226
rect 12574 544170 12642 544226
rect 12698 544170 12768 544226
rect 12448 544102 12768 544170
rect 12448 544046 12518 544102
rect 12574 544046 12642 544102
rect 12698 544046 12768 544102
rect 5418 543922 5514 543978
rect 5570 543922 5638 543978
rect 5694 543922 5762 543978
rect 5818 543922 5886 543978
rect 5942 543922 6038 543978
rect 4172 522946 4228 522956
rect 4284 530740 4340 530750
rect 4284 512484 4340 530684
rect 4284 512418 4340 512428
rect 5418 526350 6038 543922
rect 12448 543978 12768 544046
rect 12448 543922 12518 543978
rect 12574 543922 12642 543978
rect 12698 543922 12768 543978
rect 12448 543888 12768 543922
rect 43168 544350 43488 544384
rect 43168 544294 43238 544350
rect 43294 544294 43362 544350
rect 43418 544294 43488 544350
rect 43168 544226 43488 544294
rect 43168 544170 43238 544226
rect 43294 544170 43362 544226
rect 43418 544170 43488 544226
rect 43168 544102 43488 544170
rect 43168 544046 43238 544102
rect 43294 544046 43362 544102
rect 43418 544046 43488 544102
rect 43168 543978 43488 544046
rect 43168 543922 43238 543978
rect 43294 543922 43362 543978
rect 43418 543922 43488 543978
rect 43168 543888 43488 543922
rect 73888 544350 74208 544384
rect 73888 544294 73958 544350
rect 74014 544294 74082 544350
rect 74138 544294 74208 544350
rect 73888 544226 74208 544294
rect 73888 544170 73958 544226
rect 74014 544170 74082 544226
rect 74138 544170 74208 544226
rect 73888 544102 74208 544170
rect 73888 544046 73958 544102
rect 74014 544046 74082 544102
rect 74138 544046 74208 544102
rect 73888 543978 74208 544046
rect 73888 543922 73958 543978
rect 74014 543922 74082 543978
rect 74138 543922 74208 543978
rect 73888 543888 74208 543922
rect 104608 544350 104928 544384
rect 104608 544294 104678 544350
rect 104734 544294 104802 544350
rect 104858 544294 104928 544350
rect 104608 544226 104928 544294
rect 104608 544170 104678 544226
rect 104734 544170 104802 544226
rect 104858 544170 104928 544226
rect 104608 544102 104928 544170
rect 104608 544046 104678 544102
rect 104734 544046 104802 544102
rect 104858 544046 104928 544102
rect 104608 543978 104928 544046
rect 104608 543922 104678 543978
rect 104734 543922 104802 543978
rect 104858 543922 104928 543978
rect 104608 543888 104928 543922
rect 135328 544350 135648 544384
rect 135328 544294 135398 544350
rect 135454 544294 135522 544350
rect 135578 544294 135648 544350
rect 135328 544226 135648 544294
rect 135328 544170 135398 544226
rect 135454 544170 135522 544226
rect 135578 544170 135648 544226
rect 135328 544102 135648 544170
rect 135328 544046 135398 544102
rect 135454 544046 135522 544102
rect 135578 544046 135648 544102
rect 135328 543978 135648 544046
rect 135328 543922 135398 543978
rect 135454 543922 135522 543978
rect 135578 543922 135648 543978
rect 135328 543888 135648 543922
rect 166048 544350 166368 544384
rect 166048 544294 166118 544350
rect 166174 544294 166242 544350
rect 166298 544294 166368 544350
rect 166048 544226 166368 544294
rect 166048 544170 166118 544226
rect 166174 544170 166242 544226
rect 166298 544170 166368 544226
rect 166048 544102 166368 544170
rect 166048 544046 166118 544102
rect 166174 544046 166242 544102
rect 166298 544046 166368 544102
rect 166048 543978 166368 544046
rect 166048 543922 166118 543978
rect 166174 543922 166242 543978
rect 166298 543922 166368 543978
rect 166048 543888 166368 543922
rect 196768 544350 197088 544384
rect 196768 544294 196838 544350
rect 196894 544294 196962 544350
rect 197018 544294 197088 544350
rect 196768 544226 197088 544294
rect 196768 544170 196838 544226
rect 196894 544170 196962 544226
rect 197018 544170 197088 544226
rect 196768 544102 197088 544170
rect 196768 544046 196838 544102
rect 196894 544046 196962 544102
rect 197018 544046 197088 544102
rect 196768 543978 197088 544046
rect 196768 543922 196838 543978
rect 196894 543922 196962 543978
rect 197018 543922 197088 543978
rect 196768 543888 197088 543922
rect 227488 544350 227808 544384
rect 227488 544294 227558 544350
rect 227614 544294 227682 544350
rect 227738 544294 227808 544350
rect 227488 544226 227808 544294
rect 227488 544170 227558 544226
rect 227614 544170 227682 544226
rect 227738 544170 227808 544226
rect 227488 544102 227808 544170
rect 227488 544046 227558 544102
rect 227614 544046 227682 544102
rect 227738 544046 227808 544102
rect 227488 543978 227808 544046
rect 227488 543922 227558 543978
rect 227614 543922 227682 543978
rect 227738 543922 227808 543978
rect 227488 543888 227808 543922
rect 258208 544350 258528 544384
rect 258208 544294 258278 544350
rect 258334 544294 258402 544350
rect 258458 544294 258528 544350
rect 258208 544226 258528 544294
rect 258208 544170 258278 544226
rect 258334 544170 258402 544226
rect 258458 544170 258528 544226
rect 258208 544102 258528 544170
rect 258208 544046 258278 544102
rect 258334 544046 258402 544102
rect 258458 544046 258528 544102
rect 258208 543978 258528 544046
rect 258208 543922 258278 543978
rect 258334 543922 258402 543978
rect 258458 543922 258528 543978
rect 258208 543888 258528 543922
rect 288928 544350 289248 544384
rect 288928 544294 288998 544350
rect 289054 544294 289122 544350
rect 289178 544294 289248 544350
rect 288928 544226 289248 544294
rect 288928 544170 288998 544226
rect 289054 544170 289122 544226
rect 289178 544170 289248 544226
rect 288928 544102 289248 544170
rect 288928 544046 288998 544102
rect 289054 544046 289122 544102
rect 289178 544046 289248 544102
rect 288928 543978 289248 544046
rect 288928 543922 288998 543978
rect 289054 543922 289122 543978
rect 289178 543922 289248 543978
rect 288928 543888 289248 543922
rect 319648 544350 319968 544384
rect 319648 544294 319718 544350
rect 319774 544294 319842 544350
rect 319898 544294 319968 544350
rect 319648 544226 319968 544294
rect 319648 544170 319718 544226
rect 319774 544170 319842 544226
rect 319898 544170 319968 544226
rect 319648 544102 319968 544170
rect 319648 544046 319718 544102
rect 319774 544046 319842 544102
rect 319898 544046 319968 544102
rect 319648 543978 319968 544046
rect 319648 543922 319718 543978
rect 319774 543922 319842 543978
rect 319898 543922 319968 543978
rect 319648 543888 319968 543922
rect 350368 544350 350688 544384
rect 350368 544294 350438 544350
rect 350494 544294 350562 544350
rect 350618 544294 350688 544350
rect 350368 544226 350688 544294
rect 350368 544170 350438 544226
rect 350494 544170 350562 544226
rect 350618 544170 350688 544226
rect 350368 544102 350688 544170
rect 350368 544046 350438 544102
rect 350494 544046 350562 544102
rect 350618 544046 350688 544102
rect 350368 543978 350688 544046
rect 350368 543922 350438 543978
rect 350494 543922 350562 543978
rect 350618 543922 350688 543978
rect 350368 543888 350688 543922
rect 381088 544350 381408 544384
rect 381088 544294 381158 544350
rect 381214 544294 381282 544350
rect 381338 544294 381408 544350
rect 381088 544226 381408 544294
rect 381088 544170 381158 544226
rect 381214 544170 381282 544226
rect 381338 544170 381408 544226
rect 381088 544102 381408 544170
rect 381088 544046 381158 544102
rect 381214 544046 381282 544102
rect 381338 544046 381408 544102
rect 381088 543978 381408 544046
rect 381088 543922 381158 543978
rect 381214 543922 381282 543978
rect 381338 543922 381408 543978
rect 381088 543888 381408 543922
rect 411808 544350 412128 544384
rect 411808 544294 411878 544350
rect 411934 544294 412002 544350
rect 412058 544294 412128 544350
rect 411808 544226 412128 544294
rect 411808 544170 411878 544226
rect 411934 544170 412002 544226
rect 412058 544170 412128 544226
rect 411808 544102 412128 544170
rect 411808 544046 411878 544102
rect 411934 544046 412002 544102
rect 412058 544046 412128 544102
rect 411808 543978 412128 544046
rect 411808 543922 411878 543978
rect 411934 543922 412002 543978
rect 412058 543922 412128 543978
rect 411808 543888 412128 543922
rect 442528 544350 442848 544384
rect 442528 544294 442598 544350
rect 442654 544294 442722 544350
rect 442778 544294 442848 544350
rect 442528 544226 442848 544294
rect 442528 544170 442598 544226
rect 442654 544170 442722 544226
rect 442778 544170 442848 544226
rect 442528 544102 442848 544170
rect 442528 544046 442598 544102
rect 442654 544046 442722 544102
rect 442778 544046 442848 544102
rect 442528 543978 442848 544046
rect 442528 543922 442598 543978
rect 442654 543922 442722 543978
rect 442778 543922 442848 543978
rect 442528 543888 442848 543922
rect 473248 544350 473568 544384
rect 473248 544294 473318 544350
rect 473374 544294 473442 544350
rect 473498 544294 473568 544350
rect 473248 544226 473568 544294
rect 473248 544170 473318 544226
rect 473374 544170 473442 544226
rect 473498 544170 473568 544226
rect 473248 544102 473568 544170
rect 473248 544046 473318 544102
rect 473374 544046 473442 544102
rect 473498 544046 473568 544102
rect 473248 543978 473568 544046
rect 473248 543922 473318 543978
rect 473374 543922 473442 543978
rect 473498 543922 473568 543978
rect 473248 543888 473568 543922
rect 503968 544350 504288 544384
rect 503968 544294 504038 544350
rect 504094 544294 504162 544350
rect 504218 544294 504288 544350
rect 503968 544226 504288 544294
rect 503968 544170 504038 544226
rect 504094 544170 504162 544226
rect 504218 544170 504288 544226
rect 503968 544102 504288 544170
rect 503968 544046 504038 544102
rect 504094 544046 504162 544102
rect 504218 544046 504288 544102
rect 503968 543978 504288 544046
rect 503968 543922 504038 543978
rect 504094 543922 504162 543978
rect 504218 543922 504288 543978
rect 503968 543888 504288 543922
rect 534688 544350 535008 544384
rect 534688 544294 534758 544350
rect 534814 544294 534882 544350
rect 534938 544294 535008 544350
rect 534688 544226 535008 544294
rect 534688 544170 534758 544226
rect 534814 544170 534882 544226
rect 534938 544170 535008 544226
rect 534688 544102 535008 544170
rect 534688 544046 534758 544102
rect 534814 544046 534882 544102
rect 534938 544046 535008 544102
rect 534688 543978 535008 544046
rect 534688 543922 534758 543978
rect 534814 543922 534882 543978
rect 534938 543922 535008 543978
rect 534688 543888 535008 543922
rect 565408 544350 565728 544384
rect 565408 544294 565478 544350
rect 565534 544294 565602 544350
rect 565658 544294 565728 544350
rect 565408 544226 565728 544294
rect 565408 544170 565478 544226
rect 565534 544170 565602 544226
rect 565658 544170 565728 544226
rect 565408 544102 565728 544170
rect 565408 544046 565478 544102
rect 565534 544046 565602 544102
rect 565658 544046 565728 544102
rect 565408 543978 565728 544046
rect 565408 543922 565478 543978
rect 565534 543922 565602 543978
rect 565658 543922 565728 543978
rect 565408 543888 565728 543922
rect 589098 544350 589718 561922
rect 592818 550350 593438 567922
rect 592818 550294 592914 550350
rect 592970 550294 593038 550350
rect 593094 550294 593162 550350
rect 593218 550294 593286 550350
rect 593342 550294 593438 550350
rect 592818 550226 593438 550294
rect 592818 550170 592914 550226
rect 592970 550170 593038 550226
rect 593094 550170 593162 550226
rect 593218 550170 593286 550226
rect 593342 550170 593438 550226
rect 592818 550102 593438 550170
rect 592818 550046 592914 550102
rect 592970 550046 593038 550102
rect 593094 550046 593162 550102
rect 593218 550046 593286 550102
rect 593342 550046 593438 550102
rect 592818 549978 593438 550046
rect 592818 549922 592914 549978
rect 592970 549922 593038 549978
rect 593094 549922 593162 549978
rect 593218 549922 593286 549978
rect 593342 549922 593438 549978
rect 589098 544294 589194 544350
rect 589250 544294 589318 544350
rect 589374 544294 589442 544350
rect 589498 544294 589566 544350
rect 589622 544294 589718 544350
rect 589098 544226 589718 544294
rect 589098 544170 589194 544226
rect 589250 544170 589318 544226
rect 589374 544170 589442 544226
rect 589498 544170 589566 544226
rect 589622 544170 589718 544226
rect 589098 544102 589718 544170
rect 589098 544046 589194 544102
rect 589250 544046 589318 544102
rect 589374 544046 589442 544102
rect 589498 544046 589566 544102
rect 589622 544046 589718 544102
rect 589098 543978 589718 544046
rect 589098 543922 589194 543978
rect 589250 543922 589318 543978
rect 589374 543922 589442 543978
rect 589498 543922 589566 543978
rect 589622 543922 589718 543978
rect 588588 535780 588644 535790
rect 27808 532350 28128 532384
rect 27808 532294 27878 532350
rect 27934 532294 28002 532350
rect 28058 532294 28128 532350
rect 27808 532226 28128 532294
rect 27808 532170 27878 532226
rect 27934 532170 28002 532226
rect 28058 532170 28128 532226
rect 27808 532102 28128 532170
rect 27808 532046 27878 532102
rect 27934 532046 28002 532102
rect 28058 532046 28128 532102
rect 27808 531978 28128 532046
rect 27808 531922 27878 531978
rect 27934 531922 28002 531978
rect 28058 531922 28128 531978
rect 27808 531888 28128 531922
rect 58528 532350 58848 532384
rect 58528 532294 58598 532350
rect 58654 532294 58722 532350
rect 58778 532294 58848 532350
rect 58528 532226 58848 532294
rect 58528 532170 58598 532226
rect 58654 532170 58722 532226
rect 58778 532170 58848 532226
rect 58528 532102 58848 532170
rect 58528 532046 58598 532102
rect 58654 532046 58722 532102
rect 58778 532046 58848 532102
rect 58528 531978 58848 532046
rect 58528 531922 58598 531978
rect 58654 531922 58722 531978
rect 58778 531922 58848 531978
rect 58528 531888 58848 531922
rect 89248 532350 89568 532384
rect 89248 532294 89318 532350
rect 89374 532294 89442 532350
rect 89498 532294 89568 532350
rect 89248 532226 89568 532294
rect 89248 532170 89318 532226
rect 89374 532170 89442 532226
rect 89498 532170 89568 532226
rect 89248 532102 89568 532170
rect 89248 532046 89318 532102
rect 89374 532046 89442 532102
rect 89498 532046 89568 532102
rect 89248 531978 89568 532046
rect 89248 531922 89318 531978
rect 89374 531922 89442 531978
rect 89498 531922 89568 531978
rect 89248 531888 89568 531922
rect 119968 532350 120288 532384
rect 119968 532294 120038 532350
rect 120094 532294 120162 532350
rect 120218 532294 120288 532350
rect 119968 532226 120288 532294
rect 119968 532170 120038 532226
rect 120094 532170 120162 532226
rect 120218 532170 120288 532226
rect 119968 532102 120288 532170
rect 119968 532046 120038 532102
rect 120094 532046 120162 532102
rect 120218 532046 120288 532102
rect 119968 531978 120288 532046
rect 119968 531922 120038 531978
rect 120094 531922 120162 531978
rect 120218 531922 120288 531978
rect 119968 531888 120288 531922
rect 150688 532350 151008 532384
rect 150688 532294 150758 532350
rect 150814 532294 150882 532350
rect 150938 532294 151008 532350
rect 150688 532226 151008 532294
rect 150688 532170 150758 532226
rect 150814 532170 150882 532226
rect 150938 532170 151008 532226
rect 150688 532102 151008 532170
rect 150688 532046 150758 532102
rect 150814 532046 150882 532102
rect 150938 532046 151008 532102
rect 150688 531978 151008 532046
rect 150688 531922 150758 531978
rect 150814 531922 150882 531978
rect 150938 531922 151008 531978
rect 150688 531888 151008 531922
rect 181408 532350 181728 532384
rect 181408 532294 181478 532350
rect 181534 532294 181602 532350
rect 181658 532294 181728 532350
rect 181408 532226 181728 532294
rect 181408 532170 181478 532226
rect 181534 532170 181602 532226
rect 181658 532170 181728 532226
rect 181408 532102 181728 532170
rect 181408 532046 181478 532102
rect 181534 532046 181602 532102
rect 181658 532046 181728 532102
rect 181408 531978 181728 532046
rect 181408 531922 181478 531978
rect 181534 531922 181602 531978
rect 181658 531922 181728 531978
rect 181408 531888 181728 531922
rect 212128 532350 212448 532384
rect 212128 532294 212198 532350
rect 212254 532294 212322 532350
rect 212378 532294 212448 532350
rect 212128 532226 212448 532294
rect 212128 532170 212198 532226
rect 212254 532170 212322 532226
rect 212378 532170 212448 532226
rect 212128 532102 212448 532170
rect 212128 532046 212198 532102
rect 212254 532046 212322 532102
rect 212378 532046 212448 532102
rect 212128 531978 212448 532046
rect 212128 531922 212198 531978
rect 212254 531922 212322 531978
rect 212378 531922 212448 531978
rect 212128 531888 212448 531922
rect 242848 532350 243168 532384
rect 242848 532294 242918 532350
rect 242974 532294 243042 532350
rect 243098 532294 243168 532350
rect 242848 532226 243168 532294
rect 242848 532170 242918 532226
rect 242974 532170 243042 532226
rect 243098 532170 243168 532226
rect 242848 532102 243168 532170
rect 242848 532046 242918 532102
rect 242974 532046 243042 532102
rect 243098 532046 243168 532102
rect 242848 531978 243168 532046
rect 242848 531922 242918 531978
rect 242974 531922 243042 531978
rect 243098 531922 243168 531978
rect 242848 531888 243168 531922
rect 273568 532350 273888 532384
rect 273568 532294 273638 532350
rect 273694 532294 273762 532350
rect 273818 532294 273888 532350
rect 273568 532226 273888 532294
rect 273568 532170 273638 532226
rect 273694 532170 273762 532226
rect 273818 532170 273888 532226
rect 273568 532102 273888 532170
rect 273568 532046 273638 532102
rect 273694 532046 273762 532102
rect 273818 532046 273888 532102
rect 273568 531978 273888 532046
rect 273568 531922 273638 531978
rect 273694 531922 273762 531978
rect 273818 531922 273888 531978
rect 273568 531888 273888 531922
rect 304288 532350 304608 532384
rect 304288 532294 304358 532350
rect 304414 532294 304482 532350
rect 304538 532294 304608 532350
rect 304288 532226 304608 532294
rect 304288 532170 304358 532226
rect 304414 532170 304482 532226
rect 304538 532170 304608 532226
rect 304288 532102 304608 532170
rect 304288 532046 304358 532102
rect 304414 532046 304482 532102
rect 304538 532046 304608 532102
rect 304288 531978 304608 532046
rect 304288 531922 304358 531978
rect 304414 531922 304482 531978
rect 304538 531922 304608 531978
rect 304288 531888 304608 531922
rect 335008 532350 335328 532384
rect 335008 532294 335078 532350
rect 335134 532294 335202 532350
rect 335258 532294 335328 532350
rect 335008 532226 335328 532294
rect 335008 532170 335078 532226
rect 335134 532170 335202 532226
rect 335258 532170 335328 532226
rect 335008 532102 335328 532170
rect 335008 532046 335078 532102
rect 335134 532046 335202 532102
rect 335258 532046 335328 532102
rect 335008 531978 335328 532046
rect 335008 531922 335078 531978
rect 335134 531922 335202 531978
rect 335258 531922 335328 531978
rect 335008 531888 335328 531922
rect 365728 532350 366048 532384
rect 365728 532294 365798 532350
rect 365854 532294 365922 532350
rect 365978 532294 366048 532350
rect 365728 532226 366048 532294
rect 365728 532170 365798 532226
rect 365854 532170 365922 532226
rect 365978 532170 366048 532226
rect 365728 532102 366048 532170
rect 365728 532046 365798 532102
rect 365854 532046 365922 532102
rect 365978 532046 366048 532102
rect 365728 531978 366048 532046
rect 365728 531922 365798 531978
rect 365854 531922 365922 531978
rect 365978 531922 366048 531978
rect 365728 531888 366048 531922
rect 396448 532350 396768 532384
rect 396448 532294 396518 532350
rect 396574 532294 396642 532350
rect 396698 532294 396768 532350
rect 396448 532226 396768 532294
rect 396448 532170 396518 532226
rect 396574 532170 396642 532226
rect 396698 532170 396768 532226
rect 396448 532102 396768 532170
rect 396448 532046 396518 532102
rect 396574 532046 396642 532102
rect 396698 532046 396768 532102
rect 396448 531978 396768 532046
rect 396448 531922 396518 531978
rect 396574 531922 396642 531978
rect 396698 531922 396768 531978
rect 396448 531888 396768 531922
rect 427168 532350 427488 532384
rect 427168 532294 427238 532350
rect 427294 532294 427362 532350
rect 427418 532294 427488 532350
rect 427168 532226 427488 532294
rect 427168 532170 427238 532226
rect 427294 532170 427362 532226
rect 427418 532170 427488 532226
rect 427168 532102 427488 532170
rect 427168 532046 427238 532102
rect 427294 532046 427362 532102
rect 427418 532046 427488 532102
rect 427168 531978 427488 532046
rect 427168 531922 427238 531978
rect 427294 531922 427362 531978
rect 427418 531922 427488 531978
rect 427168 531888 427488 531922
rect 457888 532350 458208 532384
rect 457888 532294 457958 532350
rect 458014 532294 458082 532350
rect 458138 532294 458208 532350
rect 457888 532226 458208 532294
rect 457888 532170 457958 532226
rect 458014 532170 458082 532226
rect 458138 532170 458208 532226
rect 457888 532102 458208 532170
rect 457888 532046 457958 532102
rect 458014 532046 458082 532102
rect 458138 532046 458208 532102
rect 457888 531978 458208 532046
rect 457888 531922 457958 531978
rect 458014 531922 458082 531978
rect 458138 531922 458208 531978
rect 457888 531888 458208 531922
rect 488608 532350 488928 532384
rect 488608 532294 488678 532350
rect 488734 532294 488802 532350
rect 488858 532294 488928 532350
rect 488608 532226 488928 532294
rect 488608 532170 488678 532226
rect 488734 532170 488802 532226
rect 488858 532170 488928 532226
rect 488608 532102 488928 532170
rect 488608 532046 488678 532102
rect 488734 532046 488802 532102
rect 488858 532046 488928 532102
rect 488608 531978 488928 532046
rect 488608 531922 488678 531978
rect 488734 531922 488802 531978
rect 488858 531922 488928 531978
rect 488608 531888 488928 531922
rect 519328 532350 519648 532384
rect 519328 532294 519398 532350
rect 519454 532294 519522 532350
rect 519578 532294 519648 532350
rect 519328 532226 519648 532294
rect 519328 532170 519398 532226
rect 519454 532170 519522 532226
rect 519578 532170 519648 532226
rect 519328 532102 519648 532170
rect 519328 532046 519398 532102
rect 519454 532046 519522 532102
rect 519578 532046 519648 532102
rect 519328 531978 519648 532046
rect 519328 531922 519398 531978
rect 519454 531922 519522 531978
rect 519578 531922 519648 531978
rect 519328 531888 519648 531922
rect 550048 532350 550368 532384
rect 550048 532294 550118 532350
rect 550174 532294 550242 532350
rect 550298 532294 550368 532350
rect 550048 532226 550368 532294
rect 550048 532170 550118 532226
rect 550174 532170 550242 532226
rect 550298 532170 550368 532226
rect 550048 532102 550368 532170
rect 550048 532046 550118 532102
rect 550174 532046 550242 532102
rect 550298 532046 550368 532102
rect 550048 531978 550368 532046
rect 550048 531922 550118 531978
rect 550174 531922 550242 531978
rect 550298 531922 550368 531978
rect 550048 531888 550368 531922
rect 5418 526294 5514 526350
rect 5570 526294 5638 526350
rect 5694 526294 5762 526350
rect 5818 526294 5886 526350
rect 5942 526294 6038 526350
rect 5418 526226 6038 526294
rect 5418 526170 5514 526226
rect 5570 526170 5638 526226
rect 5694 526170 5762 526226
rect 5818 526170 5886 526226
rect 5942 526170 6038 526226
rect 5418 526102 6038 526170
rect 5418 526046 5514 526102
rect 5570 526046 5638 526102
rect 5694 526046 5762 526102
rect 5818 526046 5886 526102
rect 5942 526046 6038 526102
rect 5418 525978 6038 526046
rect 5418 525922 5514 525978
rect 5570 525922 5638 525978
rect 5694 525922 5762 525978
rect 5818 525922 5886 525978
rect 5942 525922 6038 525978
rect -956 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 -336 508350
rect -956 508226 -336 508294
rect -956 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 -336 508226
rect -956 508102 -336 508170
rect -956 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 -336 508102
rect -956 507978 -336 508046
rect -956 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 -336 507978
rect -956 490350 -336 507922
rect 5418 508350 6038 525922
rect 12448 526350 12768 526384
rect 12448 526294 12518 526350
rect 12574 526294 12642 526350
rect 12698 526294 12768 526350
rect 12448 526226 12768 526294
rect 12448 526170 12518 526226
rect 12574 526170 12642 526226
rect 12698 526170 12768 526226
rect 12448 526102 12768 526170
rect 12448 526046 12518 526102
rect 12574 526046 12642 526102
rect 12698 526046 12768 526102
rect 12448 525978 12768 526046
rect 12448 525922 12518 525978
rect 12574 525922 12642 525978
rect 12698 525922 12768 525978
rect 12448 525888 12768 525922
rect 43168 526350 43488 526384
rect 43168 526294 43238 526350
rect 43294 526294 43362 526350
rect 43418 526294 43488 526350
rect 43168 526226 43488 526294
rect 43168 526170 43238 526226
rect 43294 526170 43362 526226
rect 43418 526170 43488 526226
rect 43168 526102 43488 526170
rect 43168 526046 43238 526102
rect 43294 526046 43362 526102
rect 43418 526046 43488 526102
rect 43168 525978 43488 526046
rect 43168 525922 43238 525978
rect 43294 525922 43362 525978
rect 43418 525922 43488 525978
rect 43168 525888 43488 525922
rect 73888 526350 74208 526384
rect 73888 526294 73958 526350
rect 74014 526294 74082 526350
rect 74138 526294 74208 526350
rect 73888 526226 74208 526294
rect 73888 526170 73958 526226
rect 74014 526170 74082 526226
rect 74138 526170 74208 526226
rect 73888 526102 74208 526170
rect 73888 526046 73958 526102
rect 74014 526046 74082 526102
rect 74138 526046 74208 526102
rect 73888 525978 74208 526046
rect 73888 525922 73958 525978
rect 74014 525922 74082 525978
rect 74138 525922 74208 525978
rect 73888 525888 74208 525922
rect 104608 526350 104928 526384
rect 104608 526294 104678 526350
rect 104734 526294 104802 526350
rect 104858 526294 104928 526350
rect 104608 526226 104928 526294
rect 104608 526170 104678 526226
rect 104734 526170 104802 526226
rect 104858 526170 104928 526226
rect 104608 526102 104928 526170
rect 104608 526046 104678 526102
rect 104734 526046 104802 526102
rect 104858 526046 104928 526102
rect 104608 525978 104928 526046
rect 104608 525922 104678 525978
rect 104734 525922 104802 525978
rect 104858 525922 104928 525978
rect 104608 525888 104928 525922
rect 135328 526350 135648 526384
rect 135328 526294 135398 526350
rect 135454 526294 135522 526350
rect 135578 526294 135648 526350
rect 135328 526226 135648 526294
rect 135328 526170 135398 526226
rect 135454 526170 135522 526226
rect 135578 526170 135648 526226
rect 135328 526102 135648 526170
rect 135328 526046 135398 526102
rect 135454 526046 135522 526102
rect 135578 526046 135648 526102
rect 135328 525978 135648 526046
rect 135328 525922 135398 525978
rect 135454 525922 135522 525978
rect 135578 525922 135648 525978
rect 135328 525888 135648 525922
rect 166048 526350 166368 526384
rect 166048 526294 166118 526350
rect 166174 526294 166242 526350
rect 166298 526294 166368 526350
rect 166048 526226 166368 526294
rect 166048 526170 166118 526226
rect 166174 526170 166242 526226
rect 166298 526170 166368 526226
rect 166048 526102 166368 526170
rect 166048 526046 166118 526102
rect 166174 526046 166242 526102
rect 166298 526046 166368 526102
rect 166048 525978 166368 526046
rect 166048 525922 166118 525978
rect 166174 525922 166242 525978
rect 166298 525922 166368 525978
rect 166048 525888 166368 525922
rect 196768 526350 197088 526384
rect 196768 526294 196838 526350
rect 196894 526294 196962 526350
rect 197018 526294 197088 526350
rect 196768 526226 197088 526294
rect 196768 526170 196838 526226
rect 196894 526170 196962 526226
rect 197018 526170 197088 526226
rect 196768 526102 197088 526170
rect 196768 526046 196838 526102
rect 196894 526046 196962 526102
rect 197018 526046 197088 526102
rect 196768 525978 197088 526046
rect 196768 525922 196838 525978
rect 196894 525922 196962 525978
rect 197018 525922 197088 525978
rect 196768 525888 197088 525922
rect 227488 526350 227808 526384
rect 227488 526294 227558 526350
rect 227614 526294 227682 526350
rect 227738 526294 227808 526350
rect 227488 526226 227808 526294
rect 227488 526170 227558 526226
rect 227614 526170 227682 526226
rect 227738 526170 227808 526226
rect 227488 526102 227808 526170
rect 227488 526046 227558 526102
rect 227614 526046 227682 526102
rect 227738 526046 227808 526102
rect 227488 525978 227808 526046
rect 227488 525922 227558 525978
rect 227614 525922 227682 525978
rect 227738 525922 227808 525978
rect 227488 525888 227808 525922
rect 258208 526350 258528 526384
rect 258208 526294 258278 526350
rect 258334 526294 258402 526350
rect 258458 526294 258528 526350
rect 258208 526226 258528 526294
rect 258208 526170 258278 526226
rect 258334 526170 258402 526226
rect 258458 526170 258528 526226
rect 258208 526102 258528 526170
rect 258208 526046 258278 526102
rect 258334 526046 258402 526102
rect 258458 526046 258528 526102
rect 258208 525978 258528 526046
rect 258208 525922 258278 525978
rect 258334 525922 258402 525978
rect 258458 525922 258528 525978
rect 258208 525888 258528 525922
rect 288928 526350 289248 526384
rect 288928 526294 288998 526350
rect 289054 526294 289122 526350
rect 289178 526294 289248 526350
rect 288928 526226 289248 526294
rect 288928 526170 288998 526226
rect 289054 526170 289122 526226
rect 289178 526170 289248 526226
rect 288928 526102 289248 526170
rect 288928 526046 288998 526102
rect 289054 526046 289122 526102
rect 289178 526046 289248 526102
rect 288928 525978 289248 526046
rect 288928 525922 288998 525978
rect 289054 525922 289122 525978
rect 289178 525922 289248 525978
rect 288928 525888 289248 525922
rect 319648 526350 319968 526384
rect 319648 526294 319718 526350
rect 319774 526294 319842 526350
rect 319898 526294 319968 526350
rect 319648 526226 319968 526294
rect 319648 526170 319718 526226
rect 319774 526170 319842 526226
rect 319898 526170 319968 526226
rect 319648 526102 319968 526170
rect 319648 526046 319718 526102
rect 319774 526046 319842 526102
rect 319898 526046 319968 526102
rect 319648 525978 319968 526046
rect 319648 525922 319718 525978
rect 319774 525922 319842 525978
rect 319898 525922 319968 525978
rect 319648 525888 319968 525922
rect 350368 526350 350688 526384
rect 350368 526294 350438 526350
rect 350494 526294 350562 526350
rect 350618 526294 350688 526350
rect 350368 526226 350688 526294
rect 350368 526170 350438 526226
rect 350494 526170 350562 526226
rect 350618 526170 350688 526226
rect 350368 526102 350688 526170
rect 350368 526046 350438 526102
rect 350494 526046 350562 526102
rect 350618 526046 350688 526102
rect 350368 525978 350688 526046
rect 350368 525922 350438 525978
rect 350494 525922 350562 525978
rect 350618 525922 350688 525978
rect 350368 525888 350688 525922
rect 381088 526350 381408 526384
rect 381088 526294 381158 526350
rect 381214 526294 381282 526350
rect 381338 526294 381408 526350
rect 381088 526226 381408 526294
rect 381088 526170 381158 526226
rect 381214 526170 381282 526226
rect 381338 526170 381408 526226
rect 381088 526102 381408 526170
rect 381088 526046 381158 526102
rect 381214 526046 381282 526102
rect 381338 526046 381408 526102
rect 381088 525978 381408 526046
rect 381088 525922 381158 525978
rect 381214 525922 381282 525978
rect 381338 525922 381408 525978
rect 381088 525888 381408 525922
rect 411808 526350 412128 526384
rect 411808 526294 411878 526350
rect 411934 526294 412002 526350
rect 412058 526294 412128 526350
rect 411808 526226 412128 526294
rect 411808 526170 411878 526226
rect 411934 526170 412002 526226
rect 412058 526170 412128 526226
rect 411808 526102 412128 526170
rect 411808 526046 411878 526102
rect 411934 526046 412002 526102
rect 412058 526046 412128 526102
rect 411808 525978 412128 526046
rect 411808 525922 411878 525978
rect 411934 525922 412002 525978
rect 412058 525922 412128 525978
rect 411808 525888 412128 525922
rect 442528 526350 442848 526384
rect 442528 526294 442598 526350
rect 442654 526294 442722 526350
rect 442778 526294 442848 526350
rect 442528 526226 442848 526294
rect 442528 526170 442598 526226
rect 442654 526170 442722 526226
rect 442778 526170 442848 526226
rect 442528 526102 442848 526170
rect 442528 526046 442598 526102
rect 442654 526046 442722 526102
rect 442778 526046 442848 526102
rect 442528 525978 442848 526046
rect 442528 525922 442598 525978
rect 442654 525922 442722 525978
rect 442778 525922 442848 525978
rect 442528 525888 442848 525922
rect 473248 526350 473568 526384
rect 473248 526294 473318 526350
rect 473374 526294 473442 526350
rect 473498 526294 473568 526350
rect 473248 526226 473568 526294
rect 473248 526170 473318 526226
rect 473374 526170 473442 526226
rect 473498 526170 473568 526226
rect 473248 526102 473568 526170
rect 473248 526046 473318 526102
rect 473374 526046 473442 526102
rect 473498 526046 473568 526102
rect 473248 525978 473568 526046
rect 473248 525922 473318 525978
rect 473374 525922 473442 525978
rect 473498 525922 473568 525978
rect 473248 525888 473568 525922
rect 503968 526350 504288 526384
rect 503968 526294 504038 526350
rect 504094 526294 504162 526350
rect 504218 526294 504288 526350
rect 503968 526226 504288 526294
rect 503968 526170 504038 526226
rect 504094 526170 504162 526226
rect 504218 526170 504288 526226
rect 503968 526102 504288 526170
rect 503968 526046 504038 526102
rect 504094 526046 504162 526102
rect 504218 526046 504288 526102
rect 503968 525978 504288 526046
rect 503968 525922 504038 525978
rect 504094 525922 504162 525978
rect 504218 525922 504288 525978
rect 503968 525888 504288 525922
rect 534688 526350 535008 526384
rect 534688 526294 534758 526350
rect 534814 526294 534882 526350
rect 534938 526294 535008 526350
rect 534688 526226 535008 526294
rect 534688 526170 534758 526226
rect 534814 526170 534882 526226
rect 534938 526170 535008 526226
rect 534688 526102 535008 526170
rect 534688 526046 534758 526102
rect 534814 526046 534882 526102
rect 534938 526046 535008 526102
rect 534688 525978 535008 526046
rect 534688 525922 534758 525978
rect 534814 525922 534882 525978
rect 534938 525922 535008 525978
rect 534688 525888 535008 525922
rect 565408 526350 565728 526384
rect 565408 526294 565478 526350
rect 565534 526294 565602 526350
rect 565658 526294 565728 526350
rect 565408 526226 565728 526294
rect 565408 526170 565478 526226
rect 565534 526170 565602 526226
rect 565658 526170 565728 526226
rect 565408 526102 565728 526170
rect 565408 526046 565478 526102
rect 565534 526046 565602 526102
rect 565658 526046 565728 526102
rect 565408 525978 565728 526046
rect 565408 525922 565478 525978
rect 565534 525922 565602 525978
rect 565658 525922 565728 525978
rect 565408 525888 565728 525922
rect 588588 522564 588644 535724
rect 589098 526350 589718 543922
rect 590492 548996 590548 549006
rect 590492 533316 590548 548940
rect 590492 533250 590548 533260
rect 589098 526294 589194 526350
rect 589250 526294 589318 526350
rect 589374 526294 589442 526350
rect 589498 526294 589566 526350
rect 589622 526294 589718 526350
rect 589098 526226 589718 526294
rect 589098 526170 589194 526226
rect 589250 526170 589318 526226
rect 589374 526170 589442 526226
rect 589498 526170 589566 526226
rect 589622 526170 589718 526226
rect 589098 526102 589718 526170
rect 589098 526046 589194 526102
rect 589250 526046 589318 526102
rect 589374 526046 589442 526102
rect 589498 526046 589566 526102
rect 589622 526046 589718 526102
rect 589098 525978 589718 526046
rect 589098 525922 589194 525978
rect 589250 525922 589318 525978
rect 589374 525922 589442 525978
rect 589498 525922 589566 525978
rect 589622 525922 589718 525978
rect 588588 522498 588644 522508
rect 588812 522564 588868 522574
rect 5418 508294 5514 508350
rect 5570 508294 5638 508350
rect 5694 508294 5762 508350
rect 5818 508294 5886 508350
rect 5942 508294 6038 508350
rect 5418 508226 6038 508294
rect 5418 508170 5514 508226
rect 5570 508170 5638 508226
rect 5694 508170 5762 508226
rect 5818 508170 5886 508226
rect 5942 508170 6038 508226
rect 5418 508102 6038 508170
rect 5418 508046 5514 508102
rect 5570 508046 5638 508102
rect 5694 508046 5762 508102
rect 5818 508046 5886 508102
rect 5942 508046 6038 508102
rect 5418 507978 6038 508046
rect 5418 507922 5514 507978
rect 5570 507922 5638 507978
rect 5694 507922 5762 507978
rect 5818 507922 5886 507978
rect 5942 507922 6038 507978
rect -956 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 -336 490350
rect -956 490226 -336 490294
rect -956 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 -336 490226
rect -956 490102 -336 490170
rect -956 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 -336 490102
rect -956 489978 -336 490046
rect -956 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 -336 489978
rect -956 472350 -336 489922
rect 4172 502516 4228 502526
rect 4172 480900 4228 502460
rect 5418 490350 6038 507922
rect 6188 516628 6244 516638
rect 6188 501956 6244 516572
rect 27808 514350 28128 514384
rect 27808 514294 27878 514350
rect 27934 514294 28002 514350
rect 28058 514294 28128 514350
rect 27808 514226 28128 514294
rect 27808 514170 27878 514226
rect 27934 514170 28002 514226
rect 28058 514170 28128 514226
rect 27808 514102 28128 514170
rect 27808 514046 27878 514102
rect 27934 514046 28002 514102
rect 28058 514046 28128 514102
rect 27808 513978 28128 514046
rect 27808 513922 27878 513978
rect 27934 513922 28002 513978
rect 28058 513922 28128 513978
rect 27808 513888 28128 513922
rect 58528 514350 58848 514384
rect 58528 514294 58598 514350
rect 58654 514294 58722 514350
rect 58778 514294 58848 514350
rect 58528 514226 58848 514294
rect 58528 514170 58598 514226
rect 58654 514170 58722 514226
rect 58778 514170 58848 514226
rect 58528 514102 58848 514170
rect 58528 514046 58598 514102
rect 58654 514046 58722 514102
rect 58778 514046 58848 514102
rect 58528 513978 58848 514046
rect 58528 513922 58598 513978
rect 58654 513922 58722 513978
rect 58778 513922 58848 513978
rect 58528 513888 58848 513922
rect 89248 514350 89568 514384
rect 89248 514294 89318 514350
rect 89374 514294 89442 514350
rect 89498 514294 89568 514350
rect 89248 514226 89568 514294
rect 89248 514170 89318 514226
rect 89374 514170 89442 514226
rect 89498 514170 89568 514226
rect 89248 514102 89568 514170
rect 89248 514046 89318 514102
rect 89374 514046 89442 514102
rect 89498 514046 89568 514102
rect 89248 513978 89568 514046
rect 89248 513922 89318 513978
rect 89374 513922 89442 513978
rect 89498 513922 89568 513978
rect 89248 513888 89568 513922
rect 119968 514350 120288 514384
rect 119968 514294 120038 514350
rect 120094 514294 120162 514350
rect 120218 514294 120288 514350
rect 119968 514226 120288 514294
rect 119968 514170 120038 514226
rect 120094 514170 120162 514226
rect 120218 514170 120288 514226
rect 119968 514102 120288 514170
rect 119968 514046 120038 514102
rect 120094 514046 120162 514102
rect 120218 514046 120288 514102
rect 119968 513978 120288 514046
rect 119968 513922 120038 513978
rect 120094 513922 120162 513978
rect 120218 513922 120288 513978
rect 119968 513888 120288 513922
rect 150688 514350 151008 514384
rect 150688 514294 150758 514350
rect 150814 514294 150882 514350
rect 150938 514294 151008 514350
rect 150688 514226 151008 514294
rect 150688 514170 150758 514226
rect 150814 514170 150882 514226
rect 150938 514170 151008 514226
rect 150688 514102 151008 514170
rect 150688 514046 150758 514102
rect 150814 514046 150882 514102
rect 150938 514046 151008 514102
rect 150688 513978 151008 514046
rect 150688 513922 150758 513978
rect 150814 513922 150882 513978
rect 150938 513922 151008 513978
rect 150688 513888 151008 513922
rect 181408 514350 181728 514384
rect 181408 514294 181478 514350
rect 181534 514294 181602 514350
rect 181658 514294 181728 514350
rect 181408 514226 181728 514294
rect 181408 514170 181478 514226
rect 181534 514170 181602 514226
rect 181658 514170 181728 514226
rect 181408 514102 181728 514170
rect 181408 514046 181478 514102
rect 181534 514046 181602 514102
rect 181658 514046 181728 514102
rect 181408 513978 181728 514046
rect 181408 513922 181478 513978
rect 181534 513922 181602 513978
rect 181658 513922 181728 513978
rect 181408 513888 181728 513922
rect 212128 514350 212448 514384
rect 212128 514294 212198 514350
rect 212254 514294 212322 514350
rect 212378 514294 212448 514350
rect 212128 514226 212448 514294
rect 212128 514170 212198 514226
rect 212254 514170 212322 514226
rect 212378 514170 212448 514226
rect 212128 514102 212448 514170
rect 212128 514046 212198 514102
rect 212254 514046 212322 514102
rect 212378 514046 212448 514102
rect 212128 513978 212448 514046
rect 212128 513922 212198 513978
rect 212254 513922 212322 513978
rect 212378 513922 212448 513978
rect 212128 513888 212448 513922
rect 242848 514350 243168 514384
rect 242848 514294 242918 514350
rect 242974 514294 243042 514350
rect 243098 514294 243168 514350
rect 242848 514226 243168 514294
rect 242848 514170 242918 514226
rect 242974 514170 243042 514226
rect 243098 514170 243168 514226
rect 242848 514102 243168 514170
rect 242848 514046 242918 514102
rect 242974 514046 243042 514102
rect 243098 514046 243168 514102
rect 242848 513978 243168 514046
rect 242848 513922 242918 513978
rect 242974 513922 243042 513978
rect 243098 513922 243168 513978
rect 242848 513888 243168 513922
rect 273568 514350 273888 514384
rect 273568 514294 273638 514350
rect 273694 514294 273762 514350
rect 273818 514294 273888 514350
rect 273568 514226 273888 514294
rect 273568 514170 273638 514226
rect 273694 514170 273762 514226
rect 273818 514170 273888 514226
rect 273568 514102 273888 514170
rect 273568 514046 273638 514102
rect 273694 514046 273762 514102
rect 273818 514046 273888 514102
rect 273568 513978 273888 514046
rect 273568 513922 273638 513978
rect 273694 513922 273762 513978
rect 273818 513922 273888 513978
rect 273568 513888 273888 513922
rect 304288 514350 304608 514384
rect 304288 514294 304358 514350
rect 304414 514294 304482 514350
rect 304538 514294 304608 514350
rect 304288 514226 304608 514294
rect 304288 514170 304358 514226
rect 304414 514170 304482 514226
rect 304538 514170 304608 514226
rect 304288 514102 304608 514170
rect 304288 514046 304358 514102
rect 304414 514046 304482 514102
rect 304538 514046 304608 514102
rect 304288 513978 304608 514046
rect 304288 513922 304358 513978
rect 304414 513922 304482 513978
rect 304538 513922 304608 513978
rect 304288 513888 304608 513922
rect 335008 514350 335328 514384
rect 335008 514294 335078 514350
rect 335134 514294 335202 514350
rect 335258 514294 335328 514350
rect 335008 514226 335328 514294
rect 335008 514170 335078 514226
rect 335134 514170 335202 514226
rect 335258 514170 335328 514226
rect 335008 514102 335328 514170
rect 335008 514046 335078 514102
rect 335134 514046 335202 514102
rect 335258 514046 335328 514102
rect 335008 513978 335328 514046
rect 335008 513922 335078 513978
rect 335134 513922 335202 513978
rect 335258 513922 335328 513978
rect 335008 513888 335328 513922
rect 365728 514350 366048 514384
rect 365728 514294 365798 514350
rect 365854 514294 365922 514350
rect 365978 514294 366048 514350
rect 365728 514226 366048 514294
rect 365728 514170 365798 514226
rect 365854 514170 365922 514226
rect 365978 514170 366048 514226
rect 365728 514102 366048 514170
rect 365728 514046 365798 514102
rect 365854 514046 365922 514102
rect 365978 514046 366048 514102
rect 365728 513978 366048 514046
rect 365728 513922 365798 513978
rect 365854 513922 365922 513978
rect 365978 513922 366048 513978
rect 365728 513888 366048 513922
rect 396448 514350 396768 514384
rect 396448 514294 396518 514350
rect 396574 514294 396642 514350
rect 396698 514294 396768 514350
rect 396448 514226 396768 514294
rect 396448 514170 396518 514226
rect 396574 514170 396642 514226
rect 396698 514170 396768 514226
rect 396448 514102 396768 514170
rect 396448 514046 396518 514102
rect 396574 514046 396642 514102
rect 396698 514046 396768 514102
rect 396448 513978 396768 514046
rect 396448 513922 396518 513978
rect 396574 513922 396642 513978
rect 396698 513922 396768 513978
rect 396448 513888 396768 513922
rect 427168 514350 427488 514384
rect 427168 514294 427238 514350
rect 427294 514294 427362 514350
rect 427418 514294 427488 514350
rect 427168 514226 427488 514294
rect 427168 514170 427238 514226
rect 427294 514170 427362 514226
rect 427418 514170 427488 514226
rect 427168 514102 427488 514170
rect 427168 514046 427238 514102
rect 427294 514046 427362 514102
rect 427418 514046 427488 514102
rect 427168 513978 427488 514046
rect 427168 513922 427238 513978
rect 427294 513922 427362 513978
rect 427418 513922 427488 513978
rect 427168 513888 427488 513922
rect 457888 514350 458208 514384
rect 457888 514294 457958 514350
rect 458014 514294 458082 514350
rect 458138 514294 458208 514350
rect 457888 514226 458208 514294
rect 457888 514170 457958 514226
rect 458014 514170 458082 514226
rect 458138 514170 458208 514226
rect 457888 514102 458208 514170
rect 457888 514046 457958 514102
rect 458014 514046 458082 514102
rect 458138 514046 458208 514102
rect 457888 513978 458208 514046
rect 457888 513922 457958 513978
rect 458014 513922 458082 513978
rect 458138 513922 458208 513978
rect 457888 513888 458208 513922
rect 488608 514350 488928 514384
rect 488608 514294 488678 514350
rect 488734 514294 488802 514350
rect 488858 514294 488928 514350
rect 488608 514226 488928 514294
rect 488608 514170 488678 514226
rect 488734 514170 488802 514226
rect 488858 514170 488928 514226
rect 488608 514102 488928 514170
rect 488608 514046 488678 514102
rect 488734 514046 488802 514102
rect 488858 514046 488928 514102
rect 488608 513978 488928 514046
rect 488608 513922 488678 513978
rect 488734 513922 488802 513978
rect 488858 513922 488928 513978
rect 488608 513888 488928 513922
rect 519328 514350 519648 514384
rect 519328 514294 519398 514350
rect 519454 514294 519522 514350
rect 519578 514294 519648 514350
rect 519328 514226 519648 514294
rect 519328 514170 519398 514226
rect 519454 514170 519522 514226
rect 519578 514170 519648 514226
rect 519328 514102 519648 514170
rect 519328 514046 519398 514102
rect 519454 514046 519522 514102
rect 519578 514046 519648 514102
rect 519328 513978 519648 514046
rect 519328 513922 519398 513978
rect 519454 513922 519522 513978
rect 519578 513922 519648 513978
rect 519328 513888 519648 513922
rect 550048 514350 550368 514384
rect 550048 514294 550118 514350
rect 550174 514294 550242 514350
rect 550298 514294 550368 514350
rect 550048 514226 550368 514294
rect 550048 514170 550118 514226
rect 550174 514170 550242 514226
rect 550298 514170 550368 514226
rect 550048 514102 550368 514170
rect 550048 514046 550118 514102
rect 550174 514046 550242 514102
rect 550298 514046 550368 514102
rect 550048 513978 550368 514046
rect 550048 513922 550118 513978
rect 550174 513922 550242 513978
rect 550298 513922 550368 513978
rect 550048 513888 550368 513922
rect 588812 511812 588868 522508
rect 588812 511746 588868 511756
rect 585452 509348 585508 509358
rect 12448 508350 12768 508384
rect 12448 508294 12518 508350
rect 12574 508294 12642 508350
rect 12698 508294 12768 508350
rect 12448 508226 12768 508294
rect 12448 508170 12518 508226
rect 12574 508170 12642 508226
rect 12698 508170 12768 508226
rect 12448 508102 12768 508170
rect 12448 508046 12518 508102
rect 12574 508046 12642 508102
rect 12698 508046 12768 508102
rect 12448 507978 12768 508046
rect 12448 507922 12518 507978
rect 12574 507922 12642 507978
rect 12698 507922 12768 507978
rect 12448 507888 12768 507922
rect 43168 508350 43488 508384
rect 43168 508294 43238 508350
rect 43294 508294 43362 508350
rect 43418 508294 43488 508350
rect 43168 508226 43488 508294
rect 43168 508170 43238 508226
rect 43294 508170 43362 508226
rect 43418 508170 43488 508226
rect 43168 508102 43488 508170
rect 43168 508046 43238 508102
rect 43294 508046 43362 508102
rect 43418 508046 43488 508102
rect 43168 507978 43488 508046
rect 43168 507922 43238 507978
rect 43294 507922 43362 507978
rect 43418 507922 43488 507978
rect 43168 507888 43488 507922
rect 73888 508350 74208 508384
rect 73888 508294 73958 508350
rect 74014 508294 74082 508350
rect 74138 508294 74208 508350
rect 73888 508226 74208 508294
rect 73888 508170 73958 508226
rect 74014 508170 74082 508226
rect 74138 508170 74208 508226
rect 73888 508102 74208 508170
rect 73888 508046 73958 508102
rect 74014 508046 74082 508102
rect 74138 508046 74208 508102
rect 73888 507978 74208 508046
rect 73888 507922 73958 507978
rect 74014 507922 74082 507978
rect 74138 507922 74208 507978
rect 73888 507888 74208 507922
rect 104608 508350 104928 508384
rect 104608 508294 104678 508350
rect 104734 508294 104802 508350
rect 104858 508294 104928 508350
rect 104608 508226 104928 508294
rect 104608 508170 104678 508226
rect 104734 508170 104802 508226
rect 104858 508170 104928 508226
rect 104608 508102 104928 508170
rect 104608 508046 104678 508102
rect 104734 508046 104802 508102
rect 104858 508046 104928 508102
rect 104608 507978 104928 508046
rect 104608 507922 104678 507978
rect 104734 507922 104802 507978
rect 104858 507922 104928 507978
rect 104608 507888 104928 507922
rect 135328 508350 135648 508384
rect 135328 508294 135398 508350
rect 135454 508294 135522 508350
rect 135578 508294 135648 508350
rect 135328 508226 135648 508294
rect 135328 508170 135398 508226
rect 135454 508170 135522 508226
rect 135578 508170 135648 508226
rect 135328 508102 135648 508170
rect 135328 508046 135398 508102
rect 135454 508046 135522 508102
rect 135578 508046 135648 508102
rect 135328 507978 135648 508046
rect 135328 507922 135398 507978
rect 135454 507922 135522 507978
rect 135578 507922 135648 507978
rect 135328 507888 135648 507922
rect 166048 508350 166368 508384
rect 166048 508294 166118 508350
rect 166174 508294 166242 508350
rect 166298 508294 166368 508350
rect 166048 508226 166368 508294
rect 166048 508170 166118 508226
rect 166174 508170 166242 508226
rect 166298 508170 166368 508226
rect 166048 508102 166368 508170
rect 166048 508046 166118 508102
rect 166174 508046 166242 508102
rect 166298 508046 166368 508102
rect 166048 507978 166368 508046
rect 166048 507922 166118 507978
rect 166174 507922 166242 507978
rect 166298 507922 166368 507978
rect 166048 507888 166368 507922
rect 196768 508350 197088 508384
rect 196768 508294 196838 508350
rect 196894 508294 196962 508350
rect 197018 508294 197088 508350
rect 196768 508226 197088 508294
rect 196768 508170 196838 508226
rect 196894 508170 196962 508226
rect 197018 508170 197088 508226
rect 196768 508102 197088 508170
rect 196768 508046 196838 508102
rect 196894 508046 196962 508102
rect 197018 508046 197088 508102
rect 196768 507978 197088 508046
rect 196768 507922 196838 507978
rect 196894 507922 196962 507978
rect 197018 507922 197088 507978
rect 196768 507888 197088 507922
rect 227488 508350 227808 508384
rect 227488 508294 227558 508350
rect 227614 508294 227682 508350
rect 227738 508294 227808 508350
rect 227488 508226 227808 508294
rect 227488 508170 227558 508226
rect 227614 508170 227682 508226
rect 227738 508170 227808 508226
rect 227488 508102 227808 508170
rect 227488 508046 227558 508102
rect 227614 508046 227682 508102
rect 227738 508046 227808 508102
rect 227488 507978 227808 508046
rect 227488 507922 227558 507978
rect 227614 507922 227682 507978
rect 227738 507922 227808 507978
rect 227488 507888 227808 507922
rect 258208 508350 258528 508384
rect 258208 508294 258278 508350
rect 258334 508294 258402 508350
rect 258458 508294 258528 508350
rect 258208 508226 258528 508294
rect 258208 508170 258278 508226
rect 258334 508170 258402 508226
rect 258458 508170 258528 508226
rect 258208 508102 258528 508170
rect 258208 508046 258278 508102
rect 258334 508046 258402 508102
rect 258458 508046 258528 508102
rect 258208 507978 258528 508046
rect 258208 507922 258278 507978
rect 258334 507922 258402 507978
rect 258458 507922 258528 507978
rect 258208 507888 258528 507922
rect 288928 508350 289248 508384
rect 288928 508294 288998 508350
rect 289054 508294 289122 508350
rect 289178 508294 289248 508350
rect 288928 508226 289248 508294
rect 288928 508170 288998 508226
rect 289054 508170 289122 508226
rect 289178 508170 289248 508226
rect 288928 508102 289248 508170
rect 288928 508046 288998 508102
rect 289054 508046 289122 508102
rect 289178 508046 289248 508102
rect 288928 507978 289248 508046
rect 288928 507922 288998 507978
rect 289054 507922 289122 507978
rect 289178 507922 289248 507978
rect 288928 507888 289248 507922
rect 319648 508350 319968 508384
rect 319648 508294 319718 508350
rect 319774 508294 319842 508350
rect 319898 508294 319968 508350
rect 319648 508226 319968 508294
rect 319648 508170 319718 508226
rect 319774 508170 319842 508226
rect 319898 508170 319968 508226
rect 319648 508102 319968 508170
rect 319648 508046 319718 508102
rect 319774 508046 319842 508102
rect 319898 508046 319968 508102
rect 319648 507978 319968 508046
rect 319648 507922 319718 507978
rect 319774 507922 319842 507978
rect 319898 507922 319968 507978
rect 319648 507888 319968 507922
rect 350368 508350 350688 508384
rect 350368 508294 350438 508350
rect 350494 508294 350562 508350
rect 350618 508294 350688 508350
rect 350368 508226 350688 508294
rect 350368 508170 350438 508226
rect 350494 508170 350562 508226
rect 350618 508170 350688 508226
rect 350368 508102 350688 508170
rect 350368 508046 350438 508102
rect 350494 508046 350562 508102
rect 350618 508046 350688 508102
rect 350368 507978 350688 508046
rect 350368 507922 350438 507978
rect 350494 507922 350562 507978
rect 350618 507922 350688 507978
rect 350368 507888 350688 507922
rect 381088 508350 381408 508384
rect 381088 508294 381158 508350
rect 381214 508294 381282 508350
rect 381338 508294 381408 508350
rect 381088 508226 381408 508294
rect 381088 508170 381158 508226
rect 381214 508170 381282 508226
rect 381338 508170 381408 508226
rect 381088 508102 381408 508170
rect 381088 508046 381158 508102
rect 381214 508046 381282 508102
rect 381338 508046 381408 508102
rect 381088 507978 381408 508046
rect 381088 507922 381158 507978
rect 381214 507922 381282 507978
rect 381338 507922 381408 507978
rect 381088 507888 381408 507922
rect 411808 508350 412128 508384
rect 411808 508294 411878 508350
rect 411934 508294 412002 508350
rect 412058 508294 412128 508350
rect 411808 508226 412128 508294
rect 411808 508170 411878 508226
rect 411934 508170 412002 508226
rect 412058 508170 412128 508226
rect 411808 508102 412128 508170
rect 411808 508046 411878 508102
rect 411934 508046 412002 508102
rect 412058 508046 412128 508102
rect 411808 507978 412128 508046
rect 411808 507922 411878 507978
rect 411934 507922 412002 507978
rect 412058 507922 412128 507978
rect 411808 507888 412128 507922
rect 442528 508350 442848 508384
rect 442528 508294 442598 508350
rect 442654 508294 442722 508350
rect 442778 508294 442848 508350
rect 442528 508226 442848 508294
rect 442528 508170 442598 508226
rect 442654 508170 442722 508226
rect 442778 508170 442848 508226
rect 442528 508102 442848 508170
rect 442528 508046 442598 508102
rect 442654 508046 442722 508102
rect 442778 508046 442848 508102
rect 442528 507978 442848 508046
rect 442528 507922 442598 507978
rect 442654 507922 442722 507978
rect 442778 507922 442848 507978
rect 442528 507888 442848 507922
rect 473248 508350 473568 508384
rect 473248 508294 473318 508350
rect 473374 508294 473442 508350
rect 473498 508294 473568 508350
rect 473248 508226 473568 508294
rect 473248 508170 473318 508226
rect 473374 508170 473442 508226
rect 473498 508170 473568 508226
rect 473248 508102 473568 508170
rect 473248 508046 473318 508102
rect 473374 508046 473442 508102
rect 473498 508046 473568 508102
rect 473248 507978 473568 508046
rect 473248 507922 473318 507978
rect 473374 507922 473442 507978
rect 473498 507922 473568 507978
rect 473248 507888 473568 507922
rect 503968 508350 504288 508384
rect 503968 508294 504038 508350
rect 504094 508294 504162 508350
rect 504218 508294 504288 508350
rect 503968 508226 504288 508294
rect 503968 508170 504038 508226
rect 504094 508170 504162 508226
rect 504218 508170 504288 508226
rect 503968 508102 504288 508170
rect 503968 508046 504038 508102
rect 504094 508046 504162 508102
rect 504218 508046 504288 508102
rect 503968 507978 504288 508046
rect 503968 507922 504038 507978
rect 504094 507922 504162 507978
rect 504218 507922 504288 507978
rect 503968 507888 504288 507922
rect 534688 508350 535008 508384
rect 534688 508294 534758 508350
rect 534814 508294 534882 508350
rect 534938 508294 535008 508350
rect 534688 508226 535008 508294
rect 534688 508170 534758 508226
rect 534814 508170 534882 508226
rect 534938 508170 535008 508226
rect 534688 508102 535008 508170
rect 534688 508046 534758 508102
rect 534814 508046 534882 508102
rect 534938 508046 535008 508102
rect 534688 507978 535008 508046
rect 534688 507922 534758 507978
rect 534814 507922 534882 507978
rect 534938 507922 535008 507978
rect 534688 507888 535008 507922
rect 565408 508350 565728 508384
rect 565408 508294 565478 508350
rect 565534 508294 565602 508350
rect 565658 508294 565728 508350
rect 565408 508226 565728 508294
rect 565408 508170 565478 508226
rect 565534 508170 565602 508226
rect 565658 508170 565728 508226
rect 565408 508102 565728 508170
rect 565408 508046 565478 508102
rect 565534 508046 565602 508102
rect 565658 508046 565728 508102
rect 565408 507978 565728 508046
rect 565408 507922 565478 507978
rect 565534 507922 565602 507978
rect 565658 507922 565728 507978
rect 565408 507888 565728 507922
rect 6188 501890 6244 501900
rect 27808 496350 28128 496384
rect 27808 496294 27878 496350
rect 27934 496294 28002 496350
rect 28058 496294 28128 496350
rect 27808 496226 28128 496294
rect 27808 496170 27878 496226
rect 27934 496170 28002 496226
rect 28058 496170 28128 496226
rect 27808 496102 28128 496170
rect 27808 496046 27878 496102
rect 27934 496046 28002 496102
rect 28058 496046 28128 496102
rect 27808 495978 28128 496046
rect 27808 495922 27878 495978
rect 27934 495922 28002 495978
rect 28058 495922 28128 495978
rect 27808 495888 28128 495922
rect 58528 496350 58848 496384
rect 58528 496294 58598 496350
rect 58654 496294 58722 496350
rect 58778 496294 58848 496350
rect 58528 496226 58848 496294
rect 58528 496170 58598 496226
rect 58654 496170 58722 496226
rect 58778 496170 58848 496226
rect 58528 496102 58848 496170
rect 58528 496046 58598 496102
rect 58654 496046 58722 496102
rect 58778 496046 58848 496102
rect 58528 495978 58848 496046
rect 58528 495922 58598 495978
rect 58654 495922 58722 495978
rect 58778 495922 58848 495978
rect 58528 495888 58848 495922
rect 89248 496350 89568 496384
rect 89248 496294 89318 496350
rect 89374 496294 89442 496350
rect 89498 496294 89568 496350
rect 89248 496226 89568 496294
rect 89248 496170 89318 496226
rect 89374 496170 89442 496226
rect 89498 496170 89568 496226
rect 89248 496102 89568 496170
rect 89248 496046 89318 496102
rect 89374 496046 89442 496102
rect 89498 496046 89568 496102
rect 89248 495978 89568 496046
rect 89248 495922 89318 495978
rect 89374 495922 89442 495978
rect 89498 495922 89568 495978
rect 89248 495888 89568 495922
rect 119968 496350 120288 496384
rect 119968 496294 120038 496350
rect 120094 496294 120162 496350
rect 120218 496294 120288 496350
rect 119968 496226 120288 496294
rect 119968 496170 120038 496226
rect 120094 496170 120162 496226
rect 120218 496170 120288 496226
rect 119968 496102 120288 496170
rect 119968 496046 120038 496102
rect 120094 496046 120162 496102
rect 120218 496046 120288 496102
rect 119968 495978 120288 496046
rect 119968 495922 120038 495978
rect 120094 495922 120162 495978
rect 120218 495922 120288 495978
rect 119968 495888 120288 495922
rect 150688 496350 151008 496384
rect 150688 496294 150758 496350
rect 150814 496294 150882 496350
rect 150938 496294 151008 496350
rect 150688 496226 151008 496294
rect 150688 496170 150758 496226
rect 150814 496170 150882 496226
rect 150938 496170 151008 496226
rect 150688 496102 151008 496170
rect 150688 496046 150758 496102
rect 150814 496046 150882 496102
rect 150938 496046 151008 496102
rect 150688 495978 151008 496046
rect 150688 495922 150758 495978
rect 150814 495922 150882 495978
rect 150938 495922 151008 495978
rect 150688 495888 151008 495922
rect 181408 496350 181728 496384
rect 181408 496294 181478 496350
rect 181534 496294 181602 496350
rect 181658 496294 181728 496350
rect 181408 496226 181728 496294
rect 181408 496170 181478 496226
rect 181534 496170 181602 496226
rect 181658 496170 181728 496226
rect 181408 496102 181728 496170
rect 181408 496046 181478 496102
rect 181534 496046 181602 496102
rect 181658 496046 181728 496102
rect 181408 495978 181728 496046
rect 181408 495922 181478 495978
rect 181534 495922 181602 495978
rect 181658 495922 181728 495978
rect 181408 495888 181728 495922
rect 212128 496350 212448 496384
rect 212128 496294 212198 496350
rect 212254 496294 212322 496350
rect 212378 496294 212448 496350
rect 212128 496226 212448 496294
rect 212128 496170 212198 496226
rect 212254 496170 212322 496226
rect 212378 496170 212448 496226
rect 212128 496102 212448 496170
rect 212128 496046 212198 496102
rect 212254 496046 212322 496102
rect 212378 496046 212448 496102
rect 212128 495978 212448 496046
rect 212128 495922 212198 495978
rect 212254 495922 212322 495978
rect 212378 495922 212448 495978
rect 212128 495888 212448 495922
rect 242848 496350 243168 496384
rect 242848 496294 242918 496350
rect 242974 496294 243042 496350
rect 243098 496294 243168 496350
rect 242848 496226 243168 496294
rect 242848 496170 242918 496226
rect 242974 496170 243042 496226
rect 243098 496170 243168 496226
rect 242848 496102 243168 496170
rect 242848 496046 242918 496102
rect 242974 496046 243042 496102
rect 243098 496046 243168 496102
rect 242848 495978 243168 496046
rect 242848 495922 242918 495978
rect 242974 495922 243042 495978
rect 243098 495922 243168 495978
rect 242848 495888 243168 495922
rect 273568 496350 273888 496384
rect 273568 496294 273638 496350
rect 273694 496294 273762 496350
rect 273818 496294 273888 496350
rect 273568 496226 273888 496294
rect 273568 496170 273638 496226
rect 273694 496170 273762 496226
rect 273818 496170 273888 496226
rect 273568 496102 273888 496170
rect 273568 496046 273638 496102
rect 273694 496046 273762 496102
rect 273818 496046 273888 496102
rect 273568 495978 273888 496046
rect 273568 495922 273638 495978
rect 273694 495922 273762 495978
rect 273818 495922 273888 495978
rect 273568 495888 273888 495922
rect 304288 496350 304608 496384
rect 304288 496294 304358 496350
rect 304414 496294 304482 496350
rect 304538 496294 304608 496350
rect 304288 496226 304608 496294
rect 304288 496170 304358 496226
rect 304414 496170 304482 496226
rect 304538 496170 304608 496226
rect 304288 496102 304608 496170
rect 304288 496046 304358 496102
rect 304414 496046 304482 496102
rect 304538 496046 304608 496102
rect 304288 495978 304608 496046
rect 304288 495922 304358 495978
rect 304414 495922 304482 495978
rect 304538 495922 304608 495978
rect 304288 495888 304608 495922
rect 335008 496350 335328 496384
rect 335008 496294 335078 496350
rect 335134 496294 335202 496350
rect 335258 496294 335328 496350
rect 335008 496226 335328 496294
rect 335008 496170 335078 496226
rect 335134 496170 335202 496226
rect 335258 496170 335328 496226
rect 335008 496102 335328 496170
rect 335008 496046 335078 496102
rect 335134 496046 335202 496102
rect 335258 496046 335328 496102
rect 335008 495978 335328 496046
rect 335008 495922 335078 495978
rect 335134 495922 335202 495978
rect 335258 495922 335328 495978
rect 335008 495888 335328 495922
rect 365728 496350 366048 496384
rect 365728 496294 365798 496350
rect 365854 496294 365922 496350
rect 365978 496294 366048 496350
rect 365728 496226 366048 496294
rect 365728 496170 365798 496226
rect 365854 496170 365922 496226
rect 365978 496170 366048 496226
rect 365728 496102 366048 496170
rect 365728 496046 365798 496102
rect 365854 496046 365922 496102
rect 365978 496046 366048 496102
rect 365728 495978 366048 496046
rect 365728 495922 365798 495978
rect 365854 495922 365922 495978
rect 365978 495922 366048 495978
rect 365728 495888 366048 495922
rect 396448 496350 396768 496384
rect 396448 496294 396518 496350
rect 396574 496294 396642 496350
rect 396698 496294 396768 496350
rect 396448 496226 396768 496294
rect 396448 496170 396518 496226
rect 396574 496170 396642 496226
rect 396698 496170 396768 496226
rect 396448 496102 396768 496170
rect 396448 496046 396518 496102
rect 396574 496046 396642 496102
rect 396698 496046 396768 496102
rect 396448 495978 396768 496046
rect 396448 495922 396518 495978
rect 396574 495922 396642 495978
rect 396698 495922 396768 495978
rect 396448 495888 396768 495922
rect 427168 496350 427488 496384
rect 427168 496294 427238 496350
rect 427294 496294 427362 496350
rect 427418 496294 427488 496350
rect 427168 496226 427488 496294
rect 427168 496170 427238 496226
rect 427294 496170 427362 496226
rect 427418 496170 427488 496226
rect 427168 496102 427488 496170
rect 427168 496046 427238 496102
rect 427294 496046 427362 496102
rect 427418 496046 427488 496102
rect 427168 495978 427488 496046
rect 427168 495922 427238 495978
rect 427294 495922 427362 495978
rect 427418 495922 427488 495978
rect 427168 495888 427488 495922
rect 457888 496350 458208 496384
rect 457888 496294 457958 496350
rect 458014 496294 458082 496350
rect 458138 496294 458208 496350
rect 457888 496226 458208 496294
rect 457888 496170 457958 496226
rect 458014 496170 458082 496226
rect 458138 496170 458208 496226
rect 457888 496102 458208 496170
rect 457888 496046 457958 496102
rect 458014 496046 458082 496102
rect 458138 496046 458208 496102
rect 457888 495978 458208 496046
rect 457888 495922 457958 495978
rect 458014 495922 458082 495978
rect 458138 495922 458208 495978
rect 457888 495888 458208 495922
rect 488608 496350 488928 496384
rect 488608 496294 488678 496350
rect 488734 496294 488802 496350
rect 488858 496294 488928 496350
rect 488608 496226 488928 496294
rect 488608 496170 488678 496226
rect 488734 496170 488802 496226
rect 488858 496170 488928 496226
rect 488608 496102 488928 496170
rect 488608 496046 488678 496102
rect 488734 496046 488802 496102
rect 488858 496046 488928 496102
rect 488608 495978 488928 496046
rect 488608 495922 488678 495978
rect 488734 495922 488802 495978
rect 488858 495922 488928 495978
rect 488608 495888 488928 495922
rect 519328 496350 519648 496384
rect 519328 496294 519398 496350
rect 519454 496294 519522 496350
rect 519578 496294 519648 496350
rect 519328 496226 519648 496294
rect 519328 496170 519398 496226
rect 519454 496170 519522 496226
rect 519578 496170 519648 496226
rect 519328 496102 519648 496170
rect 519328 496046 519398 496102
rect 519454 496046 519522 496102
rect 519578 496046 519648 496102
rect 519328 495978 519648 496046
rect 519328 495922 519398 495978
rect 519454 495922 519522 495978
rect 519578 495922 519648 495978
rect 519328 495888 519648 495922
rect 550048 496350 550368 496384
rect 550048 496294 550118 496350
rect 550174 496294 550242 496350
rect 550298 496294 550368 496350
rect 550048 496226 550368 496294
rect 550048 496170 550118 496226
rect 550174 496170 550242 496226
rect 550298 496170 550368 496226
rect 550048 496102 550368 496170
rect 550048 496046 550118 496102
rect 550174 496046 550242 496102
rect 550298 496046 550368 496102
rect 550048 495978 550368 496046
rect 550048 495922 550118 495978
rect 550174 495922 550242 495978
rect 550298 495922 550368 495978
rect 550048 495888 550368 495922
rect 5418 490294 5514 490350
rect 5570 490294 5638 490350
rect 5694 490294 5762 490350
rect 5818 490294 5886 490350
rect 5942 490294 6038 490350
rect 5418 490226 6038 490294
rect 5418 490170 5514 490226
rect 5570 490170 5638 490226
rect 5694 490170 5762 490226
rect 5818 490170 5886 490226
rect 5942 490170 6038 490226
rect 5418 490102 6038 490170
rect 5418 490046 5514 490102
rect 5570 490046 5638 490102
rect 5694 490046 5762 490102
rect 5818 490046 5886 490102
rect 5942 490046 6038 490102
rect 5418 489978 6038 490046
rect 5418 489922 5514 489978
rect 5570 489922 5638 489978
rect 5694 489922 5762 489978
rect 5818 489922 5886 489978
rect 5942 489922 6038 489978
rect 4172 480834 4228 480844
rect 4284 488404 4340 488414
rect -956 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 -336 472350
rect -956 472226 -336 472294
rect -956 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 -336 472226
rect -956 472102 -336 472170
rect -956 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 -336 472102
rect -956 471978 -336 472046
rect -956 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 -336 471978
rect -956 454350 -336 471922
rect 4284 470372 4340 488348
rect 4284 470306 4340 470316
rect 5418 472350 6038 489922
rect 12448 490350 12768 490384
rect 12448 490294 12518 490350
rect 12574 490294 12642 490350
rect 12698 490294 12768 490350
rect 12448 490226 12768 490294
rect 12448 490170 12518 490226
rect 12574 490170 12642 490226
rect 12698 490170 12768 490226
rect 12448 490102 12768 490170
rect 12448 490046 12518 490102
rect 12574 490046 12642 490102
rect 12698 490046 12768 490102
rect 12448 489978 12768 490046
rect 12448 489922 12518 489978
rect 12574 489922 12642 489978
rect 12698 489922 12768 489978
rect 12448 489888 12768 489922
rect 43168 490350 43488 490384
rect 43168 490294 43238 490350
rect 43294 490294 43362 490350
rect 43418 490294 43488 490350
rect 43168 490226 43488 490294
rect 43168 490170 43238 490226
rect 43294 490170 43362 490226
rect 43418 490170 43488 490226
rect 43168 490102 43488 490170
rect 43168 490046 43238 490102
rect 43294 490046 43362 490102
rect 43418 490046 43488 490102
rect 43168 489978 43488 490046
rect 43168 489922 43238 489978
rect 43294 489922 43362 489978
rect 43418 489922 43488 489978
rect 43168 489888 43488 489922
rect 73888 490350 74208 490384
rect 73888 490294 73958 490350
rect 74014 490294 74082 490350
rect 74138 490294 74208 490350
rect 73888 490226 74208 490294
rect 73888 490170 73958 490226
rect 74014 490170 74082 490226
rect 74138 490170 74208 490226
rect 73888 490102 74208 490170
rect 73888 490046 73958 490102
rect 74014 490046 74082 490102
rect 74138 490046 74208 490102
rect 73888 489978 74208 490046
rect 73888 489922 73958 489978
rect 74014 489922 74082 489978
rect 74138 489922 74208 489978
rect 73888 489888 74208 489922
rect 104608 490350 104928 490384
rect 104608 490294 104678 490350
rect 104734 490294 104802 490350
rect 104858 490294 104928 490350
rect 104608 490226 104928 490294
rect 104608 490170 104678 490226
rect 104734 490170 104802 490226
rect 104858 490170 104928 490226
rect 104608 490102 104928 490170
rect 104608 490046 104678 490102
rect 104734 490046 104802 490102
rect 104858 490046 104928 490102
rect 104608 489978 104928 490046
rect 104608 489922 104678 489978
rect 104734 489922 104802 489978
rect 104858 489922 104928 489978
rect 104608 489888 104928 489922
rect 135328 490350 135648 490384
rect 135328 490294 135398 490350
rect 135454 490294 135522 490350
rect 135578 490294 135648 490350
rect 135328 490226 135648 490294
rect 135328 490170 135398 490226
rect 135454 490170 135522 490226
rect 135578 490170 135648 490226
rect 135328 490102 135648 490170
rect 135328 490046 135398 490102
rect 135454 490046 135522 490102
rect 135578 490046 135648 490102
rect 135328 489978 135648 490046
rect 135328 489922 135398 489978
rect 135454 489922 135522 489978
rect 135578 489922 135648 489978
rect 135328 489888 135648 489922
rect 166048 490350 166368 490384
rect 166048 490294 166118 490350
rect 166174 490294 166242 490350
rect 166298 490294 166368 490350
rect 166048 490226 166368 490294
rect 166048 490170 166118 490226
rect 166174 490170 166242 490226
rect 166298 490170 166368 490226
rect 166048 490102 166368 490170
rect 166048 490046 166118 490102
rect 166174 490046 166242 490102
rect 166298 490046 166368 490102
rect 166048 489978 166368 490046
rect 166048 489922 166118 489978
rect 166174 489922 166242 489978
rect 166298 489922 166368 489978
rect 166048 489888 166368 489922
rect 196768 490350 197088 490384
rect 196768 490294 196838 490350
rect 196894 490294 196962 490350
rect 197018 490294 197088 490350
rect 196768 490226 197088 490294
rect 196768 490170 196838 490226
rect 196894 490170 196962 490226
rect 197018 490170 197088 490226
rect 196768 490102 197088 490170
rect 196768 490046 196838 490102
rect 196894 490046 196962 490102
rect 197018 490046 197088 490102
rect 196768 489978 197088 490046
rect 196768 489922 196838 489978
rect 196894 489922 196962 489978
rect 197018 489922 197088 489978
rect 196768 489888 197088 489922
rect 227488 490350 227808 490384
rect 227488 490294 227558 490350
rect 227614 490294 227682 490350
rect 227738 490294 227808 490350
rect 227488 490226 227808 490294
rect 227488 490170 227558 490226
rect 227614 490170 227682 490226
rect 227738 490170 227808 490226
rect 227488 490102 227808 490170
rect 227488 490046 227558 490102
rect 227614 490046 227682 490102
rect 227738 490046 227808 490102
rect 227488 489978 227808 490046
rect 227488 489922 227558 489978
rect 227614 489922 227682 489978
rect 227738 489922 227808 489978
rect 227488 489888 227808 489922
rect 258208 490350 258528 490384
rect 258208 490294 258278 490350
rect 258334 490294 258402 490350
rect 258458 490294 258528 490350
rect 258208 490226 258528 490294
rect 258208 490170 258278 490226
rect 258334 490170 258402 490226
rect 258458 490170 258528 490226
rect 258208 490102 258528 490170
rect 258208 490046 258278 490102
rect 258334 490046 258402 490102
rect 258458 490046 258528 490102
rect 258208 489978 258528 490046
rect 258208 489922 258278 489978
rect 258334 489922 258402 489978
rect 258458 489922 258528 489978
rect 258208 489888 258528 489922
rect 288928 490350 289248 490384
rect 288928 490294 288998 490350
rect 289054 490294 289122 490350
rect 289178 490294 289248 490350
rect 288928 490226 289248 490294
rect 288928 490170 288998 490226
rect 289054 490170 289122 490226
rect 289178 490170 289248 490226
rect 288928 490102 289248 490170
rect 288928 490046 288998 490102
rect 289054 490046 289122 490102
rect 289178 490046 289248 490102
rect 288928 489978 289248 490046
rect 288928 489922 288998 489978
rect 289054 489922 289122 489978
rect 289178 489922 289248 489978
rect 288928 489888 289248 489922
rect 319648 490350 319968 490384
rect 319648 490294 319718 490350
rect 319774 490294 319842 490350
rect 319898 490294 319968 490350
rect 319648 490226 319968 490294
rect 319648 490170 319718 490226
rect 319774 490170 319842 490226
rect 319898 490170 319968 490226
rect 319648 490102 319968 490170
rect 319648 490046 319718 490102
rect 319774 490046 319842 490102
rect 319898 490046 319968 490102
rect 319648 489978 319968 490046
rect 319648 489922 319718 489978
rect 319774 489922 319842 489978
rect 319898 489922 319968 489978
rect 319648 489888 319968 489922
rect 350368 490350 350688 490384
rect 350368 490294 350438 490350
rect 350494 490294 350562 490350
rect 350618 490294 350688 490350
rect 350368 490226 350688 490294
rect 350368 490170 350438 490226
rect 350494 490170 350562 490226
rect 350618 490170 350688 490226
rect 350368 490102 350688 490170
rect 350368 490046 350438 490102
rect 350494 490046 350562 490102
rect 350618 490046 350688 490102
rect 350368 489978 350688 490046
rect 350368 489922 350438 489978
rect 350494 489922 350562 489978
rect 350618 489922 350688 489978
rect 350368 489888 350688 489922
rect 381088 490350 381408 490384
rect 381088 490294 381158 490350
rect 381214 490294 381282 490350
rect 381338 490294 381408 490350
rect 381088 490226 381408 490294
rect 381088 490170 381158 490226
rect 381214 490170 381282 490226
rect 381338 490170 381408 490226
rect 381088 490102 381408 490170
rect 381088 490046 381158 490102
rect 381214 490046 381282 490102
rect 381338 490046 381408 490102
rect 381088 489978 381408 490046
rect 381088 489922 381158 489978
rect 381214 489922 381282 489978
rect 381338 489922 381408 489978
rect 381088 489888 381408 489922
rect 411808 490350 412128 490384
rect 411808 490294 411878 490350
rect 411934 490294 412002 490350
rect 412058 490294 412128 490350
rect 411808 490226 412128 490294
rect 411808 490170 411878 490226
rect 411934 490170 412002 490226
rect 412058 490170 412128 490226
rect 411808 490102 412128 490170
rect 411808 490046 411878 490102
rect 411934 490046 412002 490102
rect 412058 490046 412128 490102
rect 411808 489978 412128 490046
rect 411808 489922 411878 489978
rect 411934 489922 412002 489978
rect 412058 489922 412128 489978
rect 411808 489888 412128 489922
rect 442528 490350 442848 490384
rect 442528 490294 442598 490350
rect 442654 490294 442722 490350
rect 442778 490294 442848 490350
rect 442528 490226 442848 490294
rect 442528 490170 442598 490226
rect 442654 490170 442722 490226
rect 442778 490170 442848 490226
rect 442528 490102 442848 490170
rect 442528 490046 442598 490102
rect 442654 490046 442722 490102
rect 442778 490046 442848 490102
rect 442528 489978 442848 490046
rect 442528 489922 442598 489978
rect 442654 489922 442722 489978
rect 442778 489922 442848 489978
rect 442528 489888 442848 489922
rect 473248 490350 473568 490384
rect 473248 490294 473318 490350
rect 473374 490294 473442 490350
rect 473498 490294 473568 490350
rect 473248 490226 473568 490294
rect 473248 490170 473318 490226
rect 473374 490170 473442 490226
rect 473498 490170 473568 490226
rect 473248 490102 473568 490170
rect 473248 490046 473318 490102
rect 473374 490046 473442 490102
rect 473498 490046 473568 490102
rect 473248 489978 473568 490046
rect 473248 489922 473318 489978
rect 473374 489922 473442 489978
rect 473498 489922 473568 489978
rect 473248 489888 473568 489922
rect 503968 490350 504288 490384
rect 503968 490294 504038 490350
rect 504094 490294 504162 490350
rect 504218 490294 504288 490350
rect 503968 490226 504288 490294
rect 503968 490170 504038 490226
rect 504094 490170 504162 490226
rect 504218 490170 504288 490226
rect 503968 490102 504288 490170
rect 503968 490046 504038 490102
rect 504094 490046 504162 490102
rect 504218 490046 504288 490102
rect 503968 489978 504288 490046
rect 503968 489922 504038 489978
rect 504094 489922 504162 489978
rect 504218 489922 504288 489978
rect 503968 489888 504288 489922
rect 534688 490350 535008 490384
rect 534688 490294 534758 490350
rect 534814 490294 534882 490350
rect 534938 490294 535008 490350
rect 534688 490226 535008 490294
rect 534688 490170 534758 490226
rect 534814 490170 534882 490226
rect 534938 490170 535008 490226
rect 534688 490102 535008 490170
rect 534688 490046 534758 490102
rect 534814 490046 534882 490102
rect 534938 490046 535008 490102
rect 534688 489978 535008 490046
rect 534688 489922 534758 489978
rect 534814 489922 534882 489978
rect 534938 489922 535008 489978
rect 534688 489888 535008 489922
rect 565408 490350 565728 490384
rect 565408 490294 565478 490350
rect 565534 490294 565602 490350
rect 565658 490294 565728 490350
rect 565408 490226 565728 490294
rect 585452 490308 585508 509292
rect 585452 490242 585508 490252
rect 589098 508350 589718 525922
rect 589098 508294 589194 508350
rect 589250 508294 589318 508350
rect 589374 508294 589442 508350
rect 589498 508294 589566 508350
rect 589622 508294 589718 508350
rect 589098 508226 589718 508294
rect 589098 508170 589194 508226
rect 589250 508170 589318 508226
rect 589374 508170 589442 508226
rect 589498 508170 589566 508226
rect 589622 508170 589718 508226
rect 589098 508102 589718 508170
rect 589098 508046 589194 508102
rect 589250 508046 589318 508102
rect 589374 508046 589442 508102
rect 589498 508046 589566 508102
rect 589622 508046 589718 508102
rect 589098 507978 589718 508046
rect 589098 507922 589194 507978
rect 589250 507922 589318 507978
rect 589374 507922 589442 507978
rect 589498 507922 589566 507978
rect 589622 507922 589718 507978
rect 589098 490350 589718 507922
rect 592818 532350 593438 549922
rect 592818 532294 592914 532350
rect 592970 532294 593038 532350
rect 593094 532294 593162 532350
rect 593218 532294 593286 532350
rect 593342 532294 593438 532350
rect 592818 532226 593438 532294
rect 592818 532170 592914 532226
rect 592970 532170 593038 532226
rect 593094 532170 593162 532226
rect 593218 532170 593286 532226
rect 593342 532170 593438 532226
rect 592818 532102 593438 532170
rect 592818 532046 592914 532102
rect 592970 532046 593038 532102
rect 593094 532046 593162 532102
rect 593218 532046 593286 532102
rect 593342 532046 593438 532102
rect 592818 531978 593438 532046
rect 592818 531922 592914 531978
rect 592970 531922 593038 531978
rect 593094 531922 593162 531978
rect 593218 531922 593286 531978
rect 593342 531922 593438 531978
rect 592818 514350 593438 531922
rect 592818 514294 592914 514350
rect 592970 514294 593038 514350
rect 593094 514294 593162 514350
rect 593218 514294 593286 514350
rect 593342 514294 593438 514350
rect 592818 514226 593438 514294
rect 592818 514170 592914 514226
rect 592970 514170 593038 514226
rect 593094 514170 593162 514226
rect 593218 514170 593286 514226
rect 593342 514170 593438 514226
rect 592818 514102 593438 514170
rect 592818 514046 592914 514102
rect 592970 514046 593038 514102
rect 593094 514046 593162 514102
rect 593218 514046 593286 514102
rect 593342 514046 593438 514102
rect 592818 513978 593438 514046
rect 592818 513922 592914 513978
rect 592970 513922 593038 513978
rect 593094 513922 593162 513978
rect 593218 513922 593286 513978
rect 593342 513922 593438 513978
rect 592818 496350 593438 513922
rect 592818 496294 592914 496350
rect 592970 496294 593038 496350
rect 593094 496294 593162 496350
rect 593218 496294 593286 496350
rect 593342 496294 593438 496350
rect 592818 496226 593438 496294
rect 592818 496170 592914 496226
rect 592970 496170 593038 496226
rect 593094 496170 593162 496226
rect 593218 496170 593286 496226
rect 593342 496170 593438 496226
rect 589098 490294 589194 490350
rect 589250 490294 589318 490350
rect 589374 490294 589442 490350
rect 589498 490294 589566 490350
rect 589622 490294 589718 490350
rect 565408 490170 565478 490226
rect 565534 490170 565602 490226
rect 565658 490170 565728 490226
rect 565408 490102 565728 490170
rect 565408 490046 565478 490102
rect 565534 490046 565602 490102
rect 565658 490046 565728 490102
rect 565408 489978 565728 490046
rect 565408 489922 565478 489978
rect 565534 489922 565602 489978
rect 565658 489922 565728 489978
rect 565408 489888 565728 489922
rect 589098 490226 589718 490294
rect 589098 490170 589194 490226
rect 589250 490170 589318 490226
rect 589374 490170 589442 490226
rect 589498 490170 589566 490226
rect 589622 490170 589718 490226
rect 589098 490102 589718 490170
rect 589098 490046 589194 490102
rect 589250 490046 589318 490102
rect 589374 490046 589442 490102
rect 589498 490046 589566 490102
rect 589622 490046 589718 490102
rect 589098 489978 589718 490046
rect 589098 489922 589194 489978
rect 589250 489922 589318 489978
rect 589374 489922 589442 489978
rect 589498 489922 589566 489978
rect 589622 489922 589718 489978
rect 27808 478350 28128 478384
rect 27808 478294 27878 478350
rect 27934 478294 28002 478350
rect 28058 478294 28128 478350
rect 27808 478226 28128 478294
rect 27808 478170 27878 478226
rect 27934 478170 28002 478226
rect 28058 478170 28128 478226
rect 27808 478102 28128 478170
rect 27808 478046 27878 478102
rect 27934 478046 28002 478102
rect 28058 478046 28128 478102
rect 27808 477978 28128 478046
rect 27808 477922 27878 477978
rect 27934 477922 28002 477978
rect 28058 477922 28128 477978
rect 27808 477888 28128 477922
rect 58528 478350 58848 478384
rect 58528 478294 58598 478350
rect 58654 478294 58722 478350
rect 58778 478294 58848 478350
rect 58528 478226 58848 478294
rect 58528 478170 58598 478226
rect 58654 478170 58722 478226
rect 58778 478170 58848 478226
rect 58528 478102 58848 478170
rect 58528 478046 58598 478102
rect 58654 478046 58722 478102
rect 58778 478046 58848 478102
rect 58528 477978 58848 478046
rect 58528 477922 58598 477978
rect 58654 477922 58722 477978
rect 58778 477922 58848 477978
rect 58528 477888 58848 477922
rect 89248 478350 89568 478384
rect 89248 478294 89318 478350
rect 89374 478294 89442 478350
rect 89498 478294 89568 478350
rect 89248 478226 89568 478294
rect 89248 478170 89318 478226
rect 89374 478170 89442 478226
rect 89498 478170 89568 478226
rect 89248 478102 89568 478170
rect 89248 478046 89318 478102
rect 89374 478046 89442 478102
rect 89498 478046 89568 478102
rect 89248 477978 89568 478046
rect 89248 477922 89318 477978
rect 89374 477922 89442 477978
rect 89498 477922 89568 477978
rect 89248 477888 89568 477922
rect 119968 478350 120288 478384
rect 119968 478294 120038 478350
rect 120094 478294 120162 478350
rect 120218 478294 120288 478350
rect 119968 478226 120288 478294
rect 119968 478170 120038 478226
rect 120094 478170 120162 478226
rect 120218 478170 120288 478226
rect 119968 478102 120288 478170
rect 119968 478046 120038 478102
rect 120094 478046 120162 478102
rect 120218 478046 120288 478102
rect 119968 477978 120288 478046
rect 119968 477922 120038 477978
rect 120094 477922 120162 477978
rect 120218 477922 120288 477978
rect 119968 477888 120288 477922
rect 150688 478350 151008 478384
rect 150688 478294 150758 478350
rect 150814 478294 150882 478350
rect 150938 478294 151008 478350
rect 150688 478226 151008 478294
rect 150688 478170 150758 478226
rect 150814 478170 150882 478226
rect 150938 478170 151008 478226
rect 150688 478102 151008 478170
rect 150688 478046 150758 478102
rect 150814 478046 150882 478102
rect 150938 478046 151008 478102
rect 150688 477978 151008 478046
rect 150688 477922 150758 477978
rect 150814 477922 150882 477978
rect 150938 477922 151008 477978
rect 150688 477888 151008 477922
rect 181408 478350 181728 478384
rect 181408 478294 181478 478350
rect 181534 478294 181602 478350
rect 181658 478294 181728 478350
rect 181408 478226 181728 478294
rect 181408 478170 181478 478226
rect 181534 478170 181602 478226
rect 181658 478170 181728 478226
rect 181408 478102 181728 478170
rect 181408 478046 181478 478102
rect 181534 478046 181602 478102
rect 181658 478046 181728 478102
rect 181408 477978 181728 478046
rect 181408 477922 181478 477978
rect 181534 477922 181602 477978
rect 181658 477922 181728 477978
rect 181408 477888 181728 477922
rect 212128 478350 212448 478384
rect 212128 478294 212198 478350
rect 212254 478294 212322 478350
rect 212378 478294 212448 478350
rect 212128 478226 212448 478294
rect 212128 478170 212198 478226
rect 212254 478170 212322 478226
rect 212378 478170 212448 478226
rect 212128 478102 212448 478170
rect 212128 478046 212198 478102
rect 212254 478046 212322 478102
rect 212378 478046 212448 478102
rect 212128 477978 212448 478046
rect 212128 477922 212198 477978
rect 212254 477922 212322 477978
rect 212378 477922 212448 477978
rect 212128 477888 212448 477922
rect 242848 478350 243168 478384
rect 242848 478294 242918 478350
rect 242974 478294 243042 478350
rect 243098 478294 243168 478350
rect 242848 478226 243168 478294
rect 242848 478170 242918 478226
rect 242974 478170 243042 478226
rect 243098 478170 243168 478226
rect 242848 478102 243168 478170
rect 242848 478046 242918 478102
rect 242974 478046 243042 478102
rect 243098 478046 243168 478102
rect 242848 477978 243168 478046
rect 242848 477922 242918 477978
rect 242974 477922 243042 477978
rect 243098 477922 243168 477978
rect 242848 477888 243168 477922
rect 273568 478350 273888 478384
rect 273568 478294 273638 478350
rect 273694 478294 273762 478350
rect 273818 478294 273888 478350
rect 273568 478226 273888 478294
rect 273568 478170 273638 478226
rect 273694 478170 273762 478226
rect 273818 478170 273888 478226
rect 273568 478102 273888 478170
rect 273568 478046 273638 478102
rect 273694 478046 273762 478102
rect 273818 478046 273888 478102
rect 273568 477978 273888 478046
rect 273568 477922 273638 477978
rect 273694 477922 273762 477978
rect 273818 477922 273888 477978
rect 273568 477888 273888 477922
rect 304288 478350 304608 478384
rect 304288 478294 304358 478350
rect 304414 478294 304482 478350
rect 304538 478294 304608 478350
rect 304288 478226 304608 478294
rect 304288 478170 304358 478226
rect 304414 478170 304482 478226
rect 304538 478170 304608 478226
rect 304288 478102 304608 478170
rect 304288 478046 304358 478102
rect 304414 478046 304482 478102
rect 304538 478046 304608 478102
rect 304288 477978 304608 478046
rect 304288 477922 304358 477978
rect 304414 477922 304482 477978
rect 304538 477922 304608 477978
rect 304288 477888 304608 477922
rect 335008 478350 335328 478384
rect 335008 478294 335078 478350
rect 335134 478294 335202 478350
rect 335258 478294 335328 478350
rect 335008 478226 335328 478294
rect 335008 478170 335078 478226
rect 335134 478170 335202 478226
rect 335258 478170 335328 478226
rect 335008 478102 335328 478170
rect 335008 478046 335078 478102
rect 335134 478046 335202 478102
rect 335258 478046 335328 478102
rect 335008 477978 335328 478046
rect 335008 477922 335078 477978
rect 335134 477922 335202 477978
rect 335258 477922 335328 477978
rect 335008 477888 335328 477922
rect 365728 478350 366048 478384
rect 365728 478294 365798 478350
rect 365854 478294 365922 478350
rect 365978 478294 366048 478350
rect 365728 478226 366048 478294
rect 365728 478170 365798 478226
rect 365854 478170 365922 478226
rect 365978 478170 366048 478226
rect 365728 478102 366048 478170
rect 365728 478046 365798 478102
rect 365854 478046 365922 478102
rect 365978 478046 366048 478102
rect 365728 477978 366048 478046
rect 365728 477922 365798 477978
rect 365854 477922 365922 477978
rect 365978 477922 366048 477978
rect 365728 477888 366048 477922
rect 396448 478350 396768 478384
rect 396448 478294 396518 478350
rect 396574 478294 396642 478350
rect 396698 478294 396768 478350
rect 396448 478226 396768 478294
rect 396448 478170 396518 478226
rect 396574 478170 396642 478226
rect 396698 478170 396768 478226
rect 396448 478102 396768 478170
rect 396448 478046 396518 478102
rect 396574 478046 396642 478102
rect 396698 478046 396768 478102
rect 396448 477978 396768 478046
rect 396448 477922 396518 477978
rect 396574 477922 396642 477978
rect 396698 477922 396768 477978
rect 396448 477888 396768 477922
rect 427168 478350 427488 478384
rect 427168 478294 427238 478350
rect 427294 478294 427362 478350
rect 427418 478294 427488 478350
rect 427168 478226 427488 478294
rect 427168 478170 427238 478226
rect 427294 478170 427362 478226
rect 427418 478170 427488 478226
rect 427168 478102 427488 478170
rect 427168 478046 427238 478102
rect 427294 478046 427362 478102
rect 427418 478046 427488 478102
rect 427168 477978 427488 478046
rect 427168 477922 427238 477978
rect 427294 477922 427362 477978
rect 427418 477922 427488 477978
rect 427168 477888 427488 477922
rect 457888 478350 458208 478384
rect 457888 478294 457958 478350
rect 458014 478294 458082 478350
rect 458138 478294 458208 478350
rect 457888 478226 458208 478294
rect 457888 478170 457958 478226
rect 458014 478170 458082 478226
rect 458138 478170 458208 478226
rect 457888 478102 458208 478170
rect 457888 478046 457958 478102
rect 458014 478046 458082 478102
rect 458138 478046 458208 478102
rect 457888 477978 458208 478046
rect 457888 477922 457958 477978
rect 458014 477922 458082 477978
rect 458138 477922 458208 477978
rect 457888 477888 458208 477922
rect 488608 478350 488928 478384
rect 488608 478294 488678 478350
rect 488734 478294 488802 478350
rect 488858 478294 488928 478350
rect 488608 478226 488928 478294
rect 488608 478170 488678 478226
rect 488734 478170 488802 478226
rect 488858 478170 488928 478226
rect 488608 478102 488928 478170
rect 488608 478046 488678 478102
rect 488734 478046 488802 478102
rect 488858 478046 488928 478102
rect 488608 477978 488928 478046
rect 488608 477922 488678 477978
rect 488734 477922 488802 477978
rect 488858 477922 488928 477978
rect 488608 477888 488928 477922
rect 519328 478350 519648 478384
rect 519328 478294 519398 478350
rect 519454 478294 519522 478350
rect 519578 478294 519648 478350
rect 519328 478226 519648 478294
rect 519328 478170 519398 478226
rect 519454 478170 519522 478226
rect 519578 478170 519648 478226
rect 519328 478102 519648 478170
rect 519328 478046 519398 478102
rect 519454 478046 519522 478102
rect 519578 478046 519648 478102
rect 519328 477978 519648 478046
rect 519328 477922 519398 477978
rect 519454 477922 519522 477978
rect 519578 477922 519648 477978
rect 519328 477888 519648 477922
rect 550048 478350 550368 478384
rect 550048 478294 550118 478350
rect 550174 478294 550242 478350
rect 550298 478294 550368 478350
rect 550048 478226 550368 478294
rect 550048 478170 550118 478226
rect 550174 478170 550242 478226
rect 550298 478170 550368 478226
rect 550048 478102 550368 478170
rect 550048 478046 550118 478102
rect 550174 478046 550242 478102
rect 550298 478046 550368 478102
rect 550048 477978 550368 478046
rect 550048 477922 550118 477978
rect 550174 477922 550242 477978
rect 550298 477922 550368 477978
rect 550048 477888 550368 477922
rect 5418 472294 5514 472350
rect 5570 472294 5638 472350
rect 5694 472294 5762 472350
rect 5818 472294 5886 472350
rect 5942 472294 6038 472350
rect 5418 472226 6038 472294
rect 5418 472170 5514 472226
rect 5570 472170 5638 472226
rect 5694 472170 5762 472226
rect 5818 472170 5886 472226
rect 5942 472170 6038 472226
rect 5418 472102 6038 472170
rect 5418 472046 5514 472102
rect 5570 472046 5638 472102
rect 5694 472046 5762 472102
rect 5818 472046 5886 472102
rect 5942 472046 6038 472102
rect 5418 471978 6038 472046
rect 5418 471922 5514 471978
rect 5570 471922 5638 471978
rect 5694 471922 5762 471978
rect 5818 471922 5886 471978
rect 5942 471922 6038 471978
rect -956 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 -336 454350
rect -956 454226 -336 454294
rect -956 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 -336 454226
rect -956 454102 -336 454170
rect -956 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 -336 454102
rect -956 453978 -336 454046
rect -956 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 -336 453978
rect -956 436350 -336 453922
rect 5418 454350 6038 471922
rect 6412 474292 6468 474302
rect 5418 454294 5514 454350
rect 5570 454294 5638 454350
rect 5694 454294 5762 454350
rect 5818 454294 5886 454350
rect 5942 454294 6038 454350
rect 5418 454226 6038 454294
rect 5418 454170 5514 454226
rect 5570 454170 5638 454226
rect 5694 454170 5762 454226
rect 5818 454170 5886 454226
rect 5942 454170 6038 454226
rect 5418 454102 6038 454170
rect 5418 454046 5514 454102
rect 5570 454046 5638 454102
rect 5694 454046 5762 454102
rect 5818 454046 5886 454102
rect 5942 454046 6038 454102
rect 5418 453978 6038 454046
rect 5418 453922 5514 453978
rect 5570 453922 5638 453978
rect 5694 453922 5762 453978
rect 5818 453922 5886 453978
rect 5942 453922 6038 453978
rect -956 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 -336 436350
rect -956 436226 -336 436294
rect -956 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 -336 436226
rect -956 436102 -336 436170
rect -956 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 -336 436102
rect -956 435978 -336 436046
rect -956 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 -336 435978
rect -956 418350 -336 435922
rect 4172 446068 4228 446078
rect 4172 428260 4228 446012
rect 4172 428194 4228 428204
rect 5418 436350 6038 453922
rect 6188 460180 6244 460190
rect 6188 438788 6244 460124
rect 6412 459844 6468 474236
rect 12448 472350 12768 472384
rect 12448 472294 12518 472350
rect 12574 472294 12642 472350
rect 12698 472294 12768 472350
rect 12448 472226 12768 472294
rect 12448 472170 12518 472226
rect 12574 472170 12642 472226
rect 12698 472170 12768 472226
rect 12448 472102 12768 472170
rect 12448 472046 12518 472102
rect 12574 472046 12642 472102
rect 12698 472046 12768 472102
rect 12448 471978 12768 472046
rect 12448 471922 12518 471978
rect 12574 471922 12642 471978
rect 12698 471922 12768 471978
rect 12448 471888 12768 471922
rect 43168 472350 43488 472384
rect 43168 472294 43238 472350
rect 43294 472294 43362 472350
rect 43418 472294 43488 472350
rect 43168 472226 43488 472294
rect 43168 472170 43238 472226
rect 43294 472170 43362 472226
rect 43418 472170 43488 472226
rect 43168 472102 43488 472170
rect 43168 472046 43238 472102
rect 43294 472046 43362 472102
rect 43418 472046 43488 472102
rect 43168 471978 43488 472046
rect 43168 471922 43238 471978
rect 43294 471922 43362 471978
rect 43418 471922 43488 471978
rect 43168 471888 43488 471922
rect 73888 472350 74208 472384
rect 73888 472294 73958 472350
rect 74014 472294 74082 472350
rect 74138 472294 74208 472350
rect 73888 472226 74208 472294
rect 73888 472170 73958 472226
rect 74014 472170 74082 472226
rect 74138 472170 74208 472226
rect 73888 472102 74208 472170
rect 73888 472046 73958 472102
rect 74014 472046 74082 472102
rect 74138 472046 74208 472102
rect 73888 471978 74208 472046
rect 73888 471922 73958 471978
rect 74014 471922 74082 471978
rect 74138 471922 74208 471978
rect 73888 471888 74208 471922
rect 104608 472350 104928 472384
rect 104608 472294 104678 472350
rect 104734 472294 104802 472350
rect 104858 472294 104928 472350
rect 104608 472226 104928 472294
rect 104608 472170 104678 472226
rect 104734 472170 104802 472226
rect 104858 472170 104928 472226
rect 104608 472102 104928 472170
rect 104608 472046 104678 472102
rect 104734 472046 104802 472102
rect 104858 472046 104928 472102
rect 104608 471978 104928 472046
rect 104608 471922 104678 471978
rect 104734 471922 104802 471978
rect 104858 471922 104928 471978
rect 104608 471888 104928 471922
rect 135328 472350 135648 472384
rect 135328 472294 135398 472350
rect 135454 472294 135522 472350
rect 135578 472294 135648 472350
rect 135328 472226 135648 472294
rect 135328 472170 135398 472226
rect 135454 472170 135522 472226
rect 135578 472170 135648 472226
rect 135328 472102 135648 472170
rect 135328 472046 135398 472102
rect 135454 472046 135522 472102
rect 135578 472046 135648 472102
rect 135328 471978 135648 472046
rect 135328 471922 135398 471978
rect 135454 471922 135522 471978
rect 135578 471922 135648 471978
rect 135328 471888 135648 471922
rect 166048 472350 166368 472384
rect 166048 472294 166118 472350
rect 166174 472294 166242 472350
rect 166298 472294 166368 472350
rect 166048 472226 166368 472294
rect 166048 472170 166118 472226
rect 166174 472170 166242 472226
rect 166298 472170 166368 472226
rect 166048 472102 166368 472170
rect 166048 472046 166118 472102
rect 166174 472046 166242 472102
rect 166298 472046 166368 472102
rect 166048 471978 166368 472046
rect 166048 471922 166118 471978
rect 166174 471922 166242 471978
rect 166298 471922 166368 471978
rect 166048 471888 166368 471922
rect 196768 472350 197088 472384
rect 196768 472294 196838 472350
rect 196894 472294 196962 472350
rect 197018 472294 197088 472350
rect 196768 472226 197088 472294
rect 196768 472170 196838 472226
rect 196894 472170 196962 472226
rect 197018 472170 197088 472226
rect 196768 472102 197088 472170
rect 196768 472046 196838 472102
rect 196894 472046 196962 472102
rect 197018 472046 197088 472102
rect 196768 471978 197088 472046
rect 196768 471922 196838 471978
rect 196894 471922 196962 471978
rect 197018 471922 197088 471978
rect 196768 471888 197088 471922
rect 227488 472350 227808 472384
rect 227488 472294 227558 472350
rect 227614 472294 227682 472350
rect 227738 472294 227808 472350
rect 227488 472226 227808 472294
rect 227488 472170 227558 472226
rect 227614 472170 227682 472226
rect 227738 472170 227808 472226
rect 227488 472102 227808 472170
rect 227488 472046 227558 472102
rect 227614 472046 227682 472102
rect 227738 472046 227808 472102
rect 227488 471978 227808 472046
rect 227488 471922 227558 471978
rect 227614 471922 227682 471978
rect 227738 471922 227808 471978
rect 227488 471888 227808 471922
rect 258208 472350 258528 472384
rect 258208 472294 258278 472350
rect 258334 472294 258402 472350
rect 258458 472294 258528 472350
rect 258208 472226 258528 472294
rect 258208 472170 258278 472226
rect 258334 472170 258402 472226
rect 258458 472170 258528 472226
rect 258208 472102 258528 472170
rect 258208 472046 258278 472102
rect 258334 472046 258402 472102
rect 258458 472046 258528 472102
rect 258208 471978 258528 472046
rect 258208 471922 258278 471978
rect 258334 471922 258402 471978
rect 258458 471922 258528 471978
rect 258208 471888 258528 471922
rect 288928 472350 289248 472384
rect 288928 472294 288998 472350
rect 289054 472294 289122 472350
rect 289178 472294 289248 472350
rect 288928 472226 289248 472294
rect 288928 472170 288998 472226
rect 289054 472170 289122 472226
rect 289178 472170 289248 472226
rect 288928 472102 289248 472170
rect 288928 472046 288998 472102
rect 289054 472046 289122 472102
rect 289178 472046 289248 472102
rect 288928 471978 289248 472046
rect 288928 471922 288998 471978
rect 289054 471922 289122 471978
rect 289178 471922 289248 471978
rect 288928 471888 289248 471922
rect 319648 472350 319968 472384
rect 319648 472294 319718 472350
rect 319774 472294 319842 472350
rect 319898 472294 319968 472350
rect 319648 472226 319968 472294
rect 319648 472170 319718 472226
rect 319774 472170 319842 472226
rect 319898 472170 319968 472226
rect 319648 472102 319968 472170
rect 319648 472046 319718 472102
rect 319774 472046 319842 472102
rect 319898 472046 319968 472102
rect 319648 471978 319968 472046
rect 319648 471922 319718 471978
rect 319774 471922 319842 471978
rect 319898 471922 319968 471978
rect 319648 471888 319968 471922
rect 350368 472350 350688 472384
rect 350368 472294 350438 472350
rect 350494 472294 350562 472350
rect 350618 472294 350688 472350
rect 350368 472226 350688 472294
rect 350368 472170 350438 472226
rect 350494 472170 350562 472226
rect 350618 472170 350688 472226
rect 350368 472102 350688 472170
rect 350368 472046 350438 472102
rect 350494 472046 350562 472102
rect 350618 472046 350688 472102
rect 350368 471978 350688 472046
rect 350368 471922 350438 471978
rect 350494 471922 350562 471978
rect 350618 471922 350688 471978
rect 350368 471888 350688 471922
rect 381088 472350 381408 472384
rect 381088 472294 381158 472350
rect 381214 472294 381282 472350
rect 381338 472294 381408 472350
rect 381088 472226 381408 472294
rect 381088 472170 381158 472226
rect 381214 472170 381282 472226
rect 381338 472170 381408 472226
rect 381088 472102 381408 472170
rect 381088 472046 381158 472102
rect 381214 472046 381282 472102
rect 381338 472046 381408 472102
rect 381088 471978 381408 472046
rect 381088 471922 381158 471978
rect 381214 471922 381282 471978
rect 381338 471922 381408 471978
rect 381088 471888 381408 471922
rect 411808 472350 412128 472384
rect 411808 472294 411878 472350
rect 411934 472294 412002 472350
rect 412058 472294 412128 472350
rect 411808 472226 412128 472294
rect 411808 472170 411878 472226
rect 411934 472170 412002 472226
rect 412058 472170 412128 472226
rect 411808 472102 412128 472170
rect 411808 472046 411878 472102
rect 411934 472046 412002 472102
rect 412058 472046 412128 472102
rect 411808 471978 412128 472046
rect 411808 471922 411878 471978
rect 411934 471922 412002 471978
rect 412058 471922 412128 471978
rect 411808 471888 412128 471922
rect 442528 472350 442848 472384
rect 442528 472294 442598 472350
rect 442654 472294 442722 472350
rect 442778 472294 442848 472350
rect 442528 472226 442848 472294
rect 442528 472170 442598 472226
rect 442654 472170 442722 472226
rect 442778 472170 442848 472226
rect 442528 472102 442848 472170
rect 442528 472046 442598 472102
rect 442654 472046 442722 472102
rect 442778 472046 442848 472102
rect 442528 471978 442848 472046
rect 442528 471922 442598 471978
rect 442654 471922 442722 471978
rect 442778 471922 442848 471978
rect 442528 471888 442848 471922
rect 473248 472350 473568 472384
rect 473248 472294 473318 472350
rect 473374 472294 473442 472350
rect 473498 472294 473568 472350
rect 473248 472226 473568 472294
rect 473248 472170 473318 472226
rect 473374 472170 473442 472226
rect 473498 472170 473568 472226
rect 473248 472102 473568 472170
rect 473248 472046 473318 472102
rect 473374 472046 473442 472102
rect 473498 472046 473568 472102
rect 473248 471978 473568 472046
rect 473248 471922 473318 471978
rect 473374 471922 473442 471978
rect 473498 471922 473568 471978
rect 473248 471888 473568 471922
rect 503968 472350 504288 472384
rect 503968 472294 504038 472350
rect 504094 472294 504162 472350
rect 504218 472294 504288 472350
rect 503968 472226 504288 472294
rect 503968 472170 504038 472226
rect 504094 472170 504162 472226
rect 504218 472170 504288 472226
rect 503968 472102 504288 472170
rect 503968 472046 504038 472102
rect 504094 472046 504162 472102
rect 504218 472046 504288 472102
rect 503968 471978 504288 472046
rect 503968 471922 504038 471978
rect 504094 471922 504162 471978
rect 504218 471922 504288 471978
rect 503968 471888 504288 471922
rect 534688 472350 535008 472384
rect 534688 472294 534758 472350
rect 534814 472294 534882 472350
rect 534938 472294 535008 472350
rect 534688 472226 535008 472294
rect 534688 472170 534758 472226
rect 534814 472170 534882 472226
rect 534938 472170 535008 472226
rect 534688 472102 535008 472170
rect 534688 472046 534758 472102
rect 534814 472046 534882 472102
rect 534938 472046 535008 472102
rect 534688 471978 535008 472046
rect 534688 471922 534758 471978
rect 534814 471922 534882 471978
rect 534938 471922 535008 471978
rect 534688 471888 535008 471922
rect 565408 472350 565728 472384
rect 565408 472294 565478 472350
rect 565534 472294 565602 472350
rect 565658 472294 565728 472350
rect 565408 472226 565728 472294
rect 565408 472170 565478 472226
rect 565534 472170 565602 472226
rect 565658 472170 565728 472226
rect 565408 472102 565728 472170
rect 565408 472046 565478 472102
rect 565534 472046 565602 472102
rect 565658 472046 565728 472102
rect 565408 471978 565728 472046
rect 565408 471922 565478 471978
rect 565534 471922 565602 471978
rect 565658 471922 565728 471978
rect 565408 471888 565728 471922
rect 589098 472350 589718 489922
rect 590492 496132 590548 496142
rect 590492 479556 590548 496076
rect 592818 496102 593438 496170
rect 592818 496046 592914 496102
rect 592970 496046 593038 496102
rect 593094 496046 593162 496102
rect 593218 496046 593286 496102
rect 593342 496046 593438 496102
rect 592818 495978 593438 496046
rect 592818 495922 592914 495978
rect 592970 495922 593038 495978
rect 593094 495922 593162 495978
rect 593218 495922 593286 495978
rect 593342 495922 593438 495978
rect 590492 479490 590548 479500
rect 590604 482916 590660 482926
rect 589098 472294 589194 472350
rect 589250 472294 589318 472350
rect 589374 472294 589442 472350
rect 589498 472294 589566 472350
rect 589622 472294 589718 472350
rect 589098 472226 589718 472294
rect 589098 472170 589194 472226
rect 589250 472170 589318 472226
rect 589374 472170 589442 472226
rect 589498 472170 589566 472226
rect 589622 472170 589718 472226
rect 589098 472102 589718 472170
rect 589098 472046 589194 472102
rect 589250 472046 589318 472102
rect 589374 472046 589442 472102
rect 589498 472046 589566 472102
rect 589622 472046 589718 472102
rect 589098 471978 589718 472046
rect 589098 471922 589194 471978
rect 589250 471922 589318 471978
rect 589374 471922 589442 471978
rect 589498 471922 589566 471978
rect 589622 471922 589718 471978
rect 585452 469700 585508 469710
rect 27808 460350 28128 460384
rect 27808 460294 27878 460350
rect 27934 460294 28002 460350
rect 28058 460294 28128 460350
rect 27808 460226 28128 460294
rect 27808 460170 27878 460226
rect 27934 460170 28002 460226
rect 28058 460170 28128 460226
rect 27808 460102 28128 460170
rect 27808 460046 27878 460102
rect 27934 460046 28002 460102
rect 28058 460046 28128 460102
rect 27808 459978 28128 460046
rect 27808 459922 27878 459978
rect 27934 459922 28002 459978
rect 28058 459922 28128 459978
rect 27808 459888 28128 459922
rect 58528 460350 58848 460384
rect 58528 460294 58598 460350
rect 58654 460294 58722 460350
rect 58778 460294 58848 460350
rect 58528 460226 58848 460294
rect 58528 460170 58598 460226
rect 58654 460170 58722 460226
rect 58778 460170 58848 460226
rect 58528 460102 58848 460170
rect 58528 460046 58598 460102
rect 58654 460046 58722 460102
rect 58778 460046 58848 460102
rect 58528 459978 58848 460046
rect 58528 459922 58598 459978
rect 58654 459922 58722 459978
rect 58778 459922 58848 459978
rect 58528 459888 58848 459922
rect 89248 460350 89568 460384
rect 89248 460294 89318 460350
rect 89374 460294 89442 460350
rect 89498 460294 89568 460350
rect 89248 460226 89568 460294
rect 89248 460170 89318 460226
rect 89374 460170 89442 460226
rect 89498 460170 89568 460226
rect 89248 460102 89568 460170
rect 89248 460046 89318 460102
rect 89374 460046 89442 460102
rect 89498 460046 89568 460102
rect 89248 459978 89568 460046
rect 89248 459922 89318 459978
rect 89374 459922 89442 459978
rect 89498 459922 89568 459978
rect 89248 459888 89568 459922
rect 119968 460350 120288 460384
rect 119968 460294 120038 460350
rect 120094 460294 120162 460350
rect 120218 460294 120288 460350
rect 119968 460226 120288 460294
rect 119968 460170 120038 460226
rect 120094 460170 120162 460226
rect 120218 460170 120288 460226
rect 119968 460102 120288 460170
rect 119968 460046 120038 460102
rect 120094 460046 120162 460102
rect 120218 460046 120288 460102
rect 119968 459978 120288 460046
rect 119968 459922 120038 459978
rect 120094 459922 120162 459978
rect 120218 459922 120288 459978
rect 119968 459888 120288 459922
rect 150688 460350 151008 460384
rect 150688 460294 150758 460350
rect 150814 460294 150882 460350
rect 150938 460294 151008 460350
rect 150688 460226 151008 460294
rect 150688 460170 150758 460226
rect 150814 460170 150882 460226
rect 150938 460170 151008 460226
rect 150688 460102 151008 460170
rect 150688 460046 150758 460102
rect 150814 460046 150882 460102
rect 150938 460046 151008 460102
rect 150688 459978 151008 460046
rect 150688 459922 150758 459978
rect 150814 459922 150882 459978
rect 150938 459922 151008 459978
rect 150688 459888 151008 459922
rect 181408 460350 181728 460384
rect 181408 460294 181478 460350
rect 181534 460294 181602 460350
rect 181658 460294 181728 460350
rect 181408 460226 181728 460294
rect 181408 460170 181478 460226
rect 181534 460170 181602 460226
rect 181658 460170 181728 460226
rect 181408 460102 181728 460170
rect 181408 460046 181478 460102
rect 181534 460046 181602 460102
rect 181658 460046 181728 460102
rect 181408 459978 181728 460046
rect 181408 459922 181478 459978
rect 181534 459922 181602 459978
rect 181658 459922 181728 459978
rect 181408 459888 181728 459922
rect 212128 460350 212448 460384
rect 212128 460294 212198 460350
rect 212254 460294 212322 460350
rect 212378 460294 212448 460350
rect 212128 460226 212448 460294
rect 212128 460170 212198 460226
rect 212254 460170 212322 460226
rect 212378 460170 212448 460226
rect 212128 460102 212448 460170
rect 212128 460046 212198 460102
rect 212254 460046 212322 460102
rect 212378 460046 212448 460102
rect 212128 459978 212448 460046
rect 212128 459922 212198 459978
rect 212254 459922 212322 459978
rect 212378 459922 212448 459978
rect 212128 459888 212448 459922
rect 242848 460350 243168 460384
rect 242848 460294 242918 460350
rect 242974 460294 243042 460350
rect 243098 460294 243168 460350
rect 242848 460226 243168 460294
rect 242848 460170 242918 460226
rect 242974 460170 243042 460226
rect 243098 460170 243168 460226
rect 242848 460102 243168 460170
rect 242848 460046 242918 460102
rect 242974 460046 243042 460102
rect 243098 460046 243168 460102
rect 242848 459978 243168 460046
rect 242848 459922 242918 459978
rect 242974 459922 243042 459978
rect 243098 459922 243168 459978
rect 242848 459888 243168 459922
rect 273568 460350 273888 460384
rect 273568 460294 273638 460350
rect 273694 460294 273762 460350
rect 273818 460294 273888 460350
rect 273568 460226 273888 460294
rect 273568 460170 273638 460226
rect 273694 460170 273762 460226
rect 273818 460170 273888 460226
rect 273568 460102 273888 460170
rect 273568 460046 273638 460102
rect 273694 460046 273762 460102
rect 273818 460046 273888 460102
rect 273568 459978 273888 460046
rect 273568 459922 273638 459978
rect 273694 459922 273762 459978
rect 273818 459922 273888 459978
rect 273568 459888 273888 459922
rect 304288 460350 304608 460384
rect 304288 460294 304358 460350
rect 304414 460294 304482 460350
rect 304538 460294 304608 460350
rect 304288 460226 304608 460294
rect 304288 460170 304358 460226
rect 304414 460170 304482 460226
rect 304538 460170 304608 460226
rect 304288 460102 304608 460170
rect 304288 460046 304358 460102
rect 304414 460046 304482 460102
rect 304538 460046 304608 460102
rect 304288 459978 304608 460046
rect 304288 459922 304358 459978
rect 304414 459922 304482 459978
rect 304538 459922 304608 459978
rect 304288 459888 304608 459922
rect 335008 460350 335328 460384
rect 335008 460294 335078 460350
rect 335134 460294 335202 460350
rect 335258 460294 335328 460350
rect 335008 460226 335328 460294
rect 335008 460170 335078 460226
rect 335134 460170 335202 460226
rect 335258 460170 335328 460226
rect 335008 460102 335328 460170
rect 335008 460046 335078 460102
rect 335134 460046 335202 460102
rect 335258 460046 335328 460102
rect 335008 459978 335328 460046
rect 335008 459922 335078 459978
rect 335134 459922 335202 459978
rect 335258 459922 335328 459978
rect 335008 459888 335328 459922
rect 365728 460350 366048 460384
rect 365728 460294 365798 460350
rect 365854 460294 365922 460350
rect 365978 460294 366048 460350
rect 365728 460226 366048 460294
rect 365728 460170 365798 460226
rect 365854 460170 365922 460226
rect 365978 460170 366048 460226
rect 365728 460102 366048 460170
rect 365728 460046 365798 460102
rect 365854 460046 365922 460102
rect 365978 460046 366048 460102
rect 365728 459978 366048 460046
rect 365728 459922 365798 459978
rect 365854 459922 365922 459978
rect 365978 459922 366048 459978
rect 365728 459888 366048 459922
rect 396448 460350 396768 460384
rect 396448 460294 396518 460350
rect 396574 460294 396642 460350
rect 396698 460294 396768 460350
rect 396448 460226 396768 460294
rect 396448 460170 396518 460226
rect 396574 460170 396642 460226
rect 396698 460170 396768 460226
rect 396448 460102 396768 460170
rect 396448 460046 396518 460102
rect 396574 460046 396642 460102
rect 396698 460046 396768 460102
rect 396448 459978 396768 460046
rect 396448 459922 396518 459978
rect 396574 459922 396642 459978
rect 396698 459922 396768 459978
rect 396448 459888 396768 459922
rect 427168 460350 427488 460384
rect 427168 460294 427238 460350
rect 427294 460294 427362 460350
rect 427418 460294 427488 460350
rect 427168 460226 427488 460294
rect 427168 460170 427238 460226
rect 427294 460170 427362 460226
rect 427418 460170 427488 460226
rect 427168 460102 427488 460170
rect 427168 460046 427238 460102
rect 427294 460046 427362 460102
rect 427418 460046 427488 460102
rect 427168 459978 427488 460046
rect 427168 459922 427238 459978
rect 427294 459922 427362 459978
rect 427418 459922 427488 459978
rect 427168 459888 427488 459922
rect 457888 460350 458208 460384
rect 457888 460294 457958 460350
rect 458014 460294 458082 460350
rect 458138 460294 458208 460350
rect 457888 460226 458208 460294
rect 457888 460170 457958 460226
rect 458014 460170 458082 460226
rect 458138 460170 458208 460226
rect 457888 460102 458208 460170
rect 457888 460046 457958 460102
rect 458014 460046 458082 460102
rect 458138 460046 458208 460102
rect 457888 459978 458208 460046
rect 457888 459922 457958 459978
rect 458014 459922 458082 459978
rect 458138 459922 458208 459978
rect 457888 459888 458208 459922
rect 488608 460350 488928 460384
rect 488608 460294 488678 460350
rect 488734 460294 488802 460350
rect 488858 460294 488928 460350
rect 488608 460226 488928 460294
rect 488608 460170 488678 460226
rect 488734 460170 488802 460226
rect 488858 460170 488928 460226
rect 488608 460102 488928 460170
rect 488608 460046 488678 460102
rect 488734 460046 488802 460102
rect 488858 460046 488928 460102
rect 488608 459978 488928 460046
rect 488608 459922 488678 459978
rect 488734 459922 488802 459978
rect 488858 459922 488928 459978
rect 488608 459888 488928 459922
rect 519328 460350 519648 460384
rect 519328 460294 519398 460350
rect 519454 460294 519522 460350
rect 519578 460294 519648 460350
rect 519328 460226 519648 460294
rect 519328 460170 519398 460226
rect 519454 460170 519522 460226
rect 519578 460170 519648 460226
rect 519328 460102 519648 460170
rect 519328 460046 519398 460102
rect 519454 460046 519522 460102
rect 519578 460046 519648 460102
rect 519328 459978 519648 460046
rect 519328 459922 519398 459978
rect 519454 459922 519522 459978
rect 519578 459922 519648 459978
rect 519328 459888 519648 459922
rect 550048 460350 550368 460384
rect 550048 460294 550118 460350
rect 550174 460294 550242 460350
rect 550298 460294 550368 460350
rect 550048 460226 550368 460294
rect 550048 460170 550118 460226
rect 550174 460170 550242 460226
rect 550298 460170 550368 460226
rect 550048 460102 550368 460170
rect 550048 460046 550118 460102
rect 550174 460046 550242 460102
rect 550298 460046 550368 460102
rect 550048 459978 550368 460046
rect 550048 459922 550118 459978
rect 550174 459922 550242 459978
rect 550298 459922 550368 459978
rect 550048 459888 550368 459922
rect 6412 459778 6468 459788
rect 12448 454350 12768 454384
rect 12448 454294 12518 454350
rect 12574 454294 12642 454350
rect 12698 454294 12768 454350
rect 12448 454226 12768 454294
rect 12448 454170 12518 454226
rect 12574 454170 12642 454226
rect 12698 454170 12768 454226
rect 12448 454102 12768 454170
rect 12448 454046 12518 454102
rect 12574 454046 12642 454102
rect 12698 454046 12768 454102
rect 12448 453978 12768 454046
rect 12448 453922 12518 453978
rect 12574 453922 12642 453978
rect 12698 453922 12768 453978
rect 12448 453888 12768 453922
rect 43168 454350 43488 454384
rect 43168 454294 43238 454350
rect 43294 454294 43362 454350
rect 43418 454294 43488 454350
rect 43168 454226 43488 454294
rect 43168 454170 43238 454226
rect 43294 454170 43362 454226
rect 43418 454170 43488 454226
rect 43168 454102 43488 454170
rect 43168 454046 43238 454102
rect 43294 454046 43362 454102
rect 43418 454046 43488 454102
rect 43168 453978 43488 454046
rect 43168 453922 43238 453978
rect 43294 453922 43362 453978
rect 43418 453922 43488 453978
rect 43168 453888 43488 453922
rect 73888 454350 74208 454384
rect 73888 454294 73958 454350
rect 74014 454294 74082 454350
rect 74138 454294 74208 454350
rect 73888 454226 74208 454294
rect 73888 454170 73958 454226
rect 74014 454170 74082 454226
rect 74138 454170 74208 454226
rect 73888 454102 74208 454170
rect 73888 454046 73958 454102
rect 74014 454046 74082 454102
rect 74138 454046 74208 454102
rect 73888 453978 74208 454046
rect 73888 453922 73958 453978
rect 74014 453922 74082 453978
rect 74138 453922 74208 453978
rect 73888 453888 74208 453922
rect 104608 454350 104928 454384
rect 104608 454294 104678 454350
rect 104734 454294 104802 454350
rect 104858 454294 104928 454350
rect 104608 454226 104928 454294
rect 104608 454170 104678 454226
rect 104734 454170 104802 454226
rect 104858 454170 104928 454226
rect 104608 454102 104928 454170
rect 104608 454046 104678 454102
rect 104734 454046 104802 454102
rect 104858 454046 104928 454102
rect 104608 453978 104928 454046
rect 104608 453922 104678 453978
rect 104734 453922 104802 453978
rect 104858 453922 104928 453978
rect 104608 453888 104928 453922
rect 135328 454350 135648 454384
rect 135328 454294 135398 454350
rect 135454 454294 135522 454350
rect 135578 454294 135648 454350
rect 135328 454226 135648 454294
rect 135328 454170 135398 454226
rect 135454 454170 135522 454226
rect 135578 454170 135648 454226
rect 135328 454102 135648 454170
rect 135328 454046 135398 454102
rect 135454 454046 135522 454102
rect 135578 454046 135648 454102
rect 135328 453978 135648 454046
rect 135328 453922 135398 453978
rect 135454 453922 135522 453978
rect 135578 453922 135648 453978
rect 135328 453888 135648 453922
rect 166048 454350 166368 454384
rect 166048 454294 166118 454350
rect 166174 454294 166242 454350
rect 166298 454294 166368 454350
rect 166048 454226 166368 454294
rect 166048 454170 166118 454226
rect 166174 454170 166242 454226
rect 166298 454170 166368 454226
rect 166048 454102 166368 454170
rect 166048 454046 166118 454102
rect 166174 454046 166242 454102
rect 166298 454046 166368 454102
rect 166048 453978 166368 454046
rect 166048 453922 166118 453978
rect 166174 453922 166242 453978
rect 166298 453922 166368 453978
rect 166048 453888 166368 453922
rect 196768 454350 197088 454384
rect 196768 454294 196838 454350
rect 196894 454294 196962 454350
rect 197018 454294 197088 454350
rect 196768 454226 197088 454294
rect 196768 454170 196838 454226
rect 196894 454170 196962 454226
rect 197018 454170 197088 454226
rect 196768 454102 197088 454170
rect 196768 454046 196838 454102
rect 196894 454046 196962 454102
rect 197018 454046 197088 454102
rect 196768 453978 197088 454046
rect 196768 453922 196838 453978
rect 196894 453922 196962 453978
rect 197018 453922 197088 453978
rect 196768 453888 197088 453922
rect 227488 454350 227808 454384
rect 227488 454294 227558 454350
rect 227614 454294 227682 454350
rect 227738 454294 227808 454350
rect 227488 454226 227808 454294
rect 227488 454170 227558 454226
rect 227614 454170 227682 454226
rect 227738 454170 227808 454226
rect 227488 454102 227808 454170
rect 227488 454046 227558 454102
rect 227614 454046 227682 454102
rect 227738 454046 227808 454102
rect 227488 453978 227808 454046
rect 227488 453922 227558 453978
rect 227614 453922 227682 453978
rect 227738 453922 227808 453978
rect 227488 453888 227808 453922
rect 258208 454350 258528 454384
rect 258208 454294 258278 454350
rect 258334 454294 258402 454350
rect 258458 454294 258528 454350
rect 258208 454226 258528 454294
rect 258208 454170 258278 454226
rect 258334 454170 258402 454226
rect 258458 454170 258528 454226
rect 258208 454102 258528 454170
rect 258208 454046 258278 454102
rect 258334 454046 258402 454102
rect 258458 454046 258528 454102
rect 258208 453978 258528 454046
rect 258208 453922 258278 453978
rect 258334 453922 258402 453978
rect 258458 453922 258528 453978
rect 258208 453888 258528 453922
rect 288928 454350 289248 454384
rect 288928 454294 288998 454350
rect 289054 454294 289122 454350
rect 289178 454294 289248 454350
rect 288928 454226 289248 454294
rect 288928 454170 288998 454226
rect 289054 454170 289122 454226
rect 289178 454170 289248 454226
rect 288928 454102 289248 454170
rect 288928 454046 288998 454102
rect 289054 454046 289122 454102
rect 289178 454046 289248 454102
rect 288928 453978 289248 454046
rect 288928 453922 288998 453978
rect 289054 453922 289122 453978
rect 289178 453922 289248 453978
rect 288928 453888 289248 453922
rect 319648 454350 319968 454384
rect 319648 454294 319718 454350
rect 319774 454294 319842 454350
rect 319898 454294 319968 454350
rect 319648 454226 319968 454294
rect 319648 454170 319718 454226
rect 319774 454170 319842 454226
rect 319898 454170 319968 454226
rect 319648 454102 319968 454170
rect 319648 454046 319718 454102
rect 319774 454046 319842 454102
rect 319898 454046 319968 454102
rect 319648 453978 319968 454046
rect 319648 453922 319718 453978
rect 319774 453922 319842 453978
rect 319898 453922 319968 453978
rect 319648 453888 319968 453922
rect 350368 454350 350688 454384
rect 350368 454294 350438 454350
rect 350494 454294 350562 454350
rect 350618 454294 350688 454350
rect 350368 454226 350688 454294
rect 350368 454170 350438 454226
rect 350494 454170 350562 454226
rect 350618 454170 350688 454226
rect 350368 454102 350688 454170
rect 350368 454046 350438 454102
rect 350494 454046 350562 454102
rect 350618 454046 350688 454102
rect 350368 453978 350688 454046
rect 350368 453922 350438 453978
rect 350494 453922 350562 453978
rect 350618 453922 350688 453978
rect 350368 453888 350688 453922
rect 381088 454350 381408 454384
rect 381088 454294 381158 454350
rect 381214 454294 381282 454350
rect 381338 454294 381408 454350
rect 381088 454226 381408 454294
rect 381088 454170 381158 454226
rect 381214 454170 381282 454226
rect 381338 454170 381408 454226
rect 381088 454102 381408 454170
rect 381088 454046 381158 454102
rect 381214 454046 381282 454102
rect 381338 454046 381408 454102
rect 381088 453978 381408 454046
rect 381088 453922 381158 453978
rect 381214 453922 381282 453978
rect 381338 453922 381408 453978
rect 381088 453888 381408 453922
rect 411808 454350 412128 454384
rect 411808 454294 411878 454350
rect 411934 454294 412002 454350
rect 412058 454294 412128 454350
rect 411808 454226 412128 454294
rect 411808 454170 411878 454226
rect 411934 454170 412002 454226
rect 412058 454170 412128 454226
rect 411808 454102 412128 454170
rect 411808 454046 411878 454102
rect 411934 454046 412002 454102
rect 412058 454046 412128 454102
rect 411808 453978 412128 454046
rect 411808 453922 411878 453978
rect 411934 453922 412002 453978
rect 412058 453922 412128 453978
rect 411808 453888 412128 453922
rect 442528 454350 442848 454384
rect 442528 454294 442598 454350
rect 442654 454294 442722 454350
rect 442778 454294 442848 454350
rect 442528 454226 442848 454294
rect 442528 454170 442598 454226
rect 442654 454170 442722 454226
rect 442778 454170 442848 454226
rect 442528 454102 442848 454170
rect 442528 454046 442598 454102
rect 442654 454046 442722 454102
rect 442778 454046 442848 454102
rect 442528 453978 442848 454046
rect 442528 453922 442598 453978
rect 442654 453922 442722 453978
rect 442778 453922 442848 453978
rect 442528 453888 442848 453922
rect 473248 454350 473568 454384
rect 473248 454294 473318 454350
rect 473374 454294 473442 454350
rect 473498 454294 473568 454350
rect 473248 454226 473568 454294
rect 473248 454170 473318 454226
rect 473374 454170 473442 454226
rect 473498 454170 473568 454226
rect 473248 454102 473568 454170
rect 473248 454046 473318 454102
rect 473374 454046 473442 454102
rect 473498 454046 473568 454102
rect 473248 453978 473568 454046
rect 473248 453922 473318 453978
rect 473374 453922 473442 453978
rect 473498 453922 473568 453978
rect 473248 453888 473568 453922
rect 503968 454350 504288 454384
rect 503968 454294 504038 454350
rect 504094 454294 504162 454350
rect 504218 454294 504288 454350
rect 503968 454226 504288 454294
rect 503968 454170 504038 454226
rect 504094 454170 504162 454226
rect 504218 454170 504288 454226
rect 503968 454102 504288 454170
rect 503968 454046 504038 454102
rect 504094 454046 504162 454102
rect 504218 454046 504288 454102
rect 503968 453978 504288 454046
rect 503968 453922 504038 453978
rect 504094 453922 504162 453978
rect 504218 453922 504288 453978
rect 503968 453888 504288 453922
rect 534688 454350 535008 454384
rect 534688 454294 534758 454350
rect 534814 454294 534882 454350
rect 534938 454294 535008 454350
rect 534688 454226 535008 454294
rect 534688 454170 534758 454226
rect 534814 454170 534882 454226
rect 534938 454170 535008 454226
rect 534688 454102 535008 454170
rect 534688 454046 534758 454102
rect 534814 454046 534882 454102
rect 534938 454046 535008 454102
rect 534688 453978 535008 454046
rect 534688 453922 534758 453978
rect 534814 453922 534882 453978
rect 534938 453922 535008 453978
rect 534688 453888 535008 453922
rect 565408 454350 565728 454384
rect 565408 454294 565478 454350
rect 565534 454294 565602 454350
rect 565658 454294 565728 454350
rect 565408 454226 565728 454294
rect 565408 454170 565478 454226
rect 565534 454170 565602 454226
rect 565658 454170 565728 454226
rect 565408 454102 565728 454170
rect 565408 454046 565478 454102
rect 565534 454046 565602 454102
rect 565658 454046 565728 454102
rect 565408 453978 565728 454046
rect 565408 453922 565478 453978
rect 565534 453922 565602 453978
rect 565658 453922 565728 453978
rect 565408 453888 565728 453922
rect 585452 447300 585508 469644
rect 585452 447234 585508 447244
rect 585564 456484 585620 456494
rect 27808 442350 28128 442384
rect 27808 442294 27878 442350
rect 27934 442294 28002 442350
rect 28058 442294 28128 442350
rect 27808 442226 28128 442294
rect 27808 442170 27878 442226
rect 27934 442170 28002 442226
rect 28058 442170 28128 442226
rect 27808 442102 28128 442170
rect 27808 442046 27878 442102
rect 27934 442046 28002 442102
rect 28058 442046 28128 442102
rect 27808 441978 28128 442046
rect 27808 441922 27878 441978
rect 27934 441922 28002 441978
rect 28058 441922 28128 441978
rect 27808 441888 28128 441922
rect 58528 442350 58848 442384
rect 58528 442294 58598 442350
rect 58654 442294 58722 442350
rect 58778 442294 58848 442350
rect 58528 442226 58848 442294
rect 58528 442170 58598 442226
rect 58654 442170 58722 442226
rect 58778 442170 58848 442226
rect 58528 442102 58848 442170
rect 58528 442046 58598 442102
rect 58654 442046 58722 442102
rect 58778 442046 58848 442102
rect 58528 441978 58848 442046
rect 58528 441922 58598 441978
rect 58654 441922 58722 441978
rect 58778 441922 58848 441978
rect 58528 441888 58848 441922
rect 89248 442350 89568 442384
rect 89248 442294 89318 442350
rect 89374 442294 89442 442350
rect 89498 442294 89568 442350
rect 89248 442226 89568 442294
rect 89248 442170 89318 442226
rect 89374 442170 89442 442226
rect 89498 442170 89568 442226
rect 89248 442102 89568 442170
rect 89248 442046 89318 442102
rect 89374 442046 89442 442102
rect 89498 442046 89568 442102
rect 89248 441978 89568 442046
rect 89248 441922 89318 441978
rect 89374 441922 89442 441978
rect 89498 441922 89568 441978
rect 89248 441888 89568 441922
rect 119968 442350 120288 442384
rect 119968 442294 120038 442350
rect 120094 442294 120162 442350
rect 120218 442294 120288 442350
rect 119968 442226 120288 442294
rect 119968 442170 120038 442226
rect 120094 442170 120162 442226
rect 120218 442170 120288 442226
rect 119968 442102 120288 442170
rect 119968 442046 120038 442102
rect 120094 442046 120162 442102
rect 120218 442046 120288 442102
rect 119968 441978 120288 442046
rect 119968 441922 120038 441978
rect 120094 441922 120162 441978
rect 120218 441922 120288 441978
rect 119968 441888 120288 441922
rect 150688 442350 151008 442384
rect 150688 442294 150758 442350
rect 150814 442294 150882 442350
rect 150938 442294 151008 442350
rect 150688 442226 151008 442294
rect 150688 442170 150758 442226
rect 150814 442170 150882 442226
rect 150938 442170 151008 442226
rect 150688 442102 151008 442170
rect 150688 442046 150758 442102
rect 150814 442046 150882 442102
rect 150938 442046 151008 442102
rect 150688 441978 151008 442046
rect 150688 441922 150758 441978
rect 150814 441922 150882 441978
rect 150938 441922 151008 441978
rect 150688 441888 151008 441922
rect 181408 442350 181728 442384
rect 181408 442294 181478 442350
rect 181534 442294 181602 442350
rect 181658 442294 181728 442350
rect 181408 442226 181728 442294
rect 181408 442170 181478 442226
rect 181534 442170 181602 442226
rect 181658 442170 181728 442226
rect 181408 442102 181728 442170
rect 181408 442046 181478 442102
rect 181534 442046 181602 442102
rect 181658 442046 181728 442102
rect 181408 441978 181728 442046
rect 181408 441922 181478 441978
rect 181534 441922 181602 441978
rect 181658 441922 181728 441978
rect 181408 441888 181728 441922
rect 212128 442350 212448 442384
rect 212128 442294 212198 442350
rect 212254 442294 212322 442350
rect 212378 442294 212448 442350
rect 212128 442226 212448 442294
rect 212128 442170 212198 442226
rect 212254 442170 212322 442226
rect 212378 442170 212448 442226
rect 212128 442102 212448 442170
rect 212128 442046 212198 442102
rect 212254 442046 212322 442102
rect 212378 442046 212448 442102
rect 212128 441978 212448 442046
rect 212128 441922 212198 441978
rect 212254 441922 212322 441978
rect 212378 441922 212448 441978
rect 212128 441888 212448 441922
rect 242848 442350 243168 442384
rect 242848 442294 242918 442350
rect 242974 442294 243042 442350
rect 243098 442294 243168 442350
rect 242848 442226 243168 442294
rect 242848 442170 242918 442226
rect 242974 442170 243042 442226
rect 243098 442170 243168 442226
rect 242848 442102 243168 442170
rect 242848 442046 242918 442102
rect 242974 442046 243042 442102
rect 243098 442046 243168 442102
rect 242848 441978 243168 442046
rect 242848 441922 242918 441978
rect 242974 441922 243042 441978
rect 243098 441922 243168 441978
rect 242848 441888 243168 441922
rect 273568 442350 273888 442384
rect 273568 442294 273638 442350
rect 273694 442294 273762 442350
rect 273818 442294 273888 442350
rect 273568 442226 273888 442294
rect 273568 442170 273638 442226
rect 273694 442170 273762 442226
rect 273818 442170 273888 442226
rect 273568 442102 273888 442170
rect 273568 442046 273638 442102
rect 273694 442046 273762 442102
rect 273818 442046 273888 442102
rect 273568 441978 273888 442046
rect 273568 441922 273638 441978
rect 273694 441922 273762 441978
rect 273818 441922 273888 441978
rect 273568 441888 273888 441922
rect 304288 442350 304608 442384
rect 304288 442294 304358 442350
rect 304414 442294 304482 442350
rect 304538 442294 304608 442350
rect 304288 442226 304608 442294
rect 304288 442170 304358 442226
rect 304414 442170 304482 442226
rect 304538 442170 304608 442226
rect 304288 442102 304608 442170
rect 304288 442046 304358 442102
rect 304414 442046 304482 442102
rect 304538 442046 304608 442102
rect 304288 441978 304608 442046
rect 304288 441922 304358 441978
rect 304414 441922 304482 441978
rect 304538 441922 304608 441978
rect 304288 441888 304608 441922
rect 335008 442350 335328 442384
rect 335008 442294 335078 442350
rect 335134 442294 335202 442350
rect 335258 442294 335328 442350
rect 335008 442226 335328 442294
rect 335008 442170 335078 442226
rect 335134 442170 335202 442226
rect 335258 442170 335328 442226
rect 335008 442102 335328 442170
rect 335008 442046 335078 442102
rect 335134 442046 335202 442102
rect 335258 442046 335328 442102
rect 335008 441978 335328 442046
rect 335008 441922 335078 441978
rect 335134 441922 335202 441978
rect 335258 441922 335328 441978
rect 335008 441888 335328 441922
rect 365728 442350 366048 442384
rect 365728 442294 365798 442350
rect 365854 442294 365922 442350
rect 365978 442294 366048 442350
rect 365728 442226 366048 442294
rect 365728 442170 365798 442226
rect 365854 442170 365922 442226
rect 365978 442170 366048 442226
rect 365728 442102 366048 442170
rect 365728 442046 365798 442102
rect 365854 442046 365922 442102
rect 365978 442046 366048 442102
rect 365728 441978 366048 442046
rect 365728 441922 365798 441978
rect 365854 441922 365922 441978
rect 365978 441922 366048 441978
rect 365728 441888 366048 441922
rect 396448 442350 396768 442384
rect 396448 442294 396518 442350
rect 396574 442294 396642 442350
rect 396698 442294 396768 442350
rect 396448 442226 396768 442294
rect 396448 442170 396518 442226
rect 396574 442170 396642 442226
rect 396698 442170 396768 442226
rect 396448 442102 396768 442170
rect 396448 442046 396518 442102
rect 396574 442046 396642 442102
rect 396698 442046 396768 442102
rect 396448 441978 396768 442046
rect 396448 441922 396518 441978
rect 396574 441922 396642 441978
rect 396698 441922 396768 441978
rect 396448 441888 396768 441922
rect 427168 442350 427488 442384
rect 427168 442294 427238 442350
rect 427294 442294 427362 442350
rect 427418 442294 427488 442350
rect 427168 442226 427488 442294
rect 427168 442170 427238 442226
rect 427294 442170 427362 442226
rect 427418 442170 427488 442226
rect 427168 442102 427488 442170
rect 427168 442046 427238 442102
rect 427294 442046 427362 442102
rect 427418 442046 427488 442102
rect 427168 441978 427488 442046
rect 427168 441922 427238 441978
rect 427294 441922 427362 441978
rect 427418 441922 427488 441978
rect 427168 441888 427488 441922
rect 457888 442350 458208 442384
rect 457888 442294 457958 442350
rect 458014 442294 458082 442350
rect 458138 442294 458208 442350
rect 457888 442226 458208 442294
rect 457888 442170 457958 442226
rect 458014 442170 458082 442226
rect 458138 442170 458208 442226
rect 457888 442102 458208 442170
rect 457888 442046 457958 442102
rect 458014 442046 458082 442102
rect 458138 442046 458208 442102
rect 457888 441978 458208 442046
rect 457888 441922 457958 441978
rect 458014 441922 458082 441978
rect 458138 441922 458208 441978
rect 457888 441888 458208 441922
rect 488608 442350 488928 442384
rect 488608 442294 488678 442350
rect 488734 442294 488802 442350
rect 488858 442294 488928 442350
rect 488608 442226 488928 442294
rect 488608 442170 488678 442226
rect 488734 442170 488802 442226
rect 488858 442170 488928 442226
rect 488608 442102 488928 442170
rect 488608 442046 488678 442102
rect 488734 442046 488802 442102
rect 488858 442046 488928 442102
rect 488608 441978 488928 442046
rect 488608 441922 488678 441978
rect 488734 441922 488802 441978
rect 488858 441922 488928 441978
rect 488608 441888 488928 441922
rect 519328 442350 519648 442384
rect 519328 442294 519398 442350
rect 519454 442294 519522 442350
rect 519578 442294 519648 442350
rect 519328 442226 519648 442294
rect 519328 442170 519398 442226
rect 519454 442170 519522 442226
rect 519578 442170 519648 442226
rect 519328 442102 519648 442170
rect 519328 442046 519398 442102
rect 519454 442046 519522 442102
rect 519578 442046 519648 442102
rect 519328 441978 519648 442046
rect 519328 441922 519398 441978
rect 519454 441922 519522 441978
rect 519578 441922 519648 441978
rect 519328 441888 519648 441922
rect 550048 442350 550368 442384
rect 550048 442294 550118 442350
rect 550174 442294 550242 442350
rect 550298 442294 550368 442350
rect 550048 442226 550368 442294
rect 550048 442170 550118 442226
rect 550174 442170 550242 442226
rect 550298 442170 550368 442226
rect 550048 442102 550368 442170
rect 550048 442046 550118 442102
rect 550174 442046 550242 442102
rect 550298 442046 550368 442102
rect 550048 441978 550368 442046
rect 550048 441922 550118 441978
rect 550174 441922 550242 441978
rect 550298 441922 550368 441978
rect 550048 441888 550368 441922
rect 6188 438722 6244 438732
rect 585564 436548 585620 456428
rect 585564 436482 585620 436492
rect 589098 454350 589718 471922
rect 590604 468804 590660 482860
rect 590604 468738 590660 468748
rect 592818 478350 593438 495922
rect 592818 478294 592914 478350
rect 592970 478294 593038 478350
rect 593094 478294 593162 478350
rect 593218 478294 593286 478350
rect 593342 478294 593438 478350
rect 592818 478226 593438 478294
rect 592818 478170 592914 478226
rect 592970 478170 593038 478226
rect 593094 478170 593162 478226
rect 593218 478170 593286 478226
rect 593342 478170 593438 478226
rect 592818 478102 593438 478170
rect 592818 478046 592914 478102
rect 592970 478046 593038 478102
rect 593094 478046 593162 478102
rect 593218 478046 593286 478102
rect 593342 478046 593438 478102
rect 592818 477978 593438 478046
rect 592818 477922 592914 477978
rect 592970 477922 593038 477978
rect 593094 477922 593162 477978
rect 593218 477922 593286 477978
rect 593342 477922 593438 477978
rect 589098 454294 589194 454350
rect 589250 454294 589318 454350
rect 589374 454294 589442 454350
rect 589498 454294 589566 454350
rect 589622 454294 589718 454350
rect 589098 454226 589718 454294
rect 589098 454170 589194 454226
rect 589250 454170 589318 454226
rect 589374 454170 589442 454226
rect 589498 454170 589566 454226
rect 589622 454170 589718 454226
rect 589098 454102 589718 454170
rect 589098 454046 589194 454102
rect 589250 454046 589318 454102
rect 589374 454046 589442 454102
rect 589498 454046 589566 454102
rect 589622 454046 589718 454102
rect 589098 453978 589718 454046
rect 589098 453922 589194 453978
rect 589250 453922 589318 453978
rect 589374 453922 589442 453978
rect 589498 453922 589566 453978
rect 589622 453922 589718 453978
rect 5418 436294 5514 436350
rect 5570 436294 5638 436350
rect 5694 436294 5762 436350
rect 5818 436294 5886 436350
rect 5942 436294 6038 436350
rect 5418 436226 6038 436294
rect 5418 436170 5514 436226
rect 5570 436170 5638 436226
rect 5694 436170 5762 436226
rect 5818 436170 5886 436226
rect 5942 436170 6038 436226
rect 5418 436102 6038 436170
rect 5418 436046 5514 436102
rect 5570 436046 5638 436102
rect 5694 436046 5762 436102
rect 5818 436046 5886 436102
rect 5942 436046 6038 436102
rect 5418 435978 6038 436046
rect 5418 435922 5514 435978
rect 5570 435922 5638 435978
rect 5694 435922 5762 435978
rect 5818 435922 5886 435978
rect 5942 435922 6038 435978
rect -956 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 -336 418350
rect -956 418226 -336 418294
rect -956 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 -336 418226
rect -956 418102 -336 418170
rect -956 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 -336 418102
rect -956 417978 -336 418046
rect -956 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 -336 417978
rect -956 400350 -336 417922
rect 5418 418350 6038 435922
rect 12448 436350 12768 436384
rect 12448 436294 12518 436350
rect 12574 436294 12642 436350
rect 12698 436294 12768 436350
rect 12448 436226 12768 436294
rect 12448 436170 12518 436226
rect 12574 436170 12642 436226
rect 12698 436170 12768 436226
rect 12448 436102 12768 436170
rect 12448 436046 12518 436102
rect 12574 436046 12642 436102
rect 12698 436046 12768 436102
rect 12448 435978 12768 436046
rect 12448 435922 12518 435978
rect 12574 435922 12642 435978
rect 12698 435922 12768 435978
rect 12448 435888 12768 435922
rect 43168 436350 43488 436384
rect 43168 436294 43238 436350
rect 43294 436294 43362 436350
rect 43418 436294 43488 436350
rect 43168 436226 43488 436294
rect 43168 436170 43238 436226
rect 43294 436170 43362 436226
rect 43418 436170 43488 436226
rect 43168 436102 43488 436170
rect 43168 436046 43238 436102
rect 43294 436046 43362 436102
rect 43418 436046 43488 436102
rect 43168 435978 43488 436046
rect 43168 435922 43238 435978
rect 43294 435922 43362 435978
rect 43418 435922 43488 435978
rect 43168 435888 43488 435922
rect 73888 436350 74208 436384
rect 73888 436294 73958 436350
rect 74014 436294 74082 436350
rect 74138 436294 74208 436350
rect 73888 436226 74208 436294
rect 73888 436170 73958 436226
rect 74014 436170 74082 436226
rect 74138 436170 74208 436226
rect 73888 436102 74208 436170
rect 73888 436046 73958 436102
rect 74014 436046 74082 436102
rect 74138 436046 74208 436102
rect 73888 435978 74208 436046
rect 73888 435922 73958 435978
rect 74014 435922 74082 435978
rect 74138 435922 74208 435978
rect 73888 435888 74208 435922
rect 104608 436350 104928 436384
rect 104608 436294 104678 436350
rect 104734 436294 104802 436350
rect 104858 436294 104928 436350
rect 104608 436226 104928 436294
rect 104608 436170 104678 436226
rect 104734 436170 104802 436226
rect 104858 436170 104928 436226
rect 104608 436102 104928 436170
rect 104608 436046 104678 436102
rect 104734 436046 104802 436102
rect 104858 436046 104928 436102
rect 104608 435978 104928 436046
rect 104608 435922 104678 435978
rect 104734 435922 104802 435978
rect 104858 435922 104928 435978
rect 104608 435888 104928 435922
rect 135328 436350 135648 436384
rect 135328 436294 135398 436350
rect 135454 436294 135522 436350
rect 135578 436294 135648 436350
rect 135328 436226 135648 436294
rect 135328 436170 135398 436226
rect 135454 436170 135522 436226
rect 135578 436170 135648 436226
rect 135328 436102 135648 436170
rect 135328 436046 135398 436102
rect 135454 436046 135522 436102
rect 135578 436046 135648 436102
rect 135328 435978 135648 436046
rect 135328 435922 135398 435978
rect 135454 435922 135522 435978
rect 135578 435922 135648 435978
rect 135328 435888 135648 435922
rect 166048 436350 166368 436384
rect 166048 436294 166118 436350
rect 166174 436294 166242 436350
rect 166298 436294 166368 436350
rect 166048 436226 166368 436294
rect 166048 436170 166118 436226
rect 166174 436170 166242 436226
rect 166298 436170 166368 436226
rect 166048 436102 166368 436170
rect 166048 436046 166118 436102
rect 166174 436046 166242 436102
rect 166298 436046 166368 436102
rect 166048 435978 166368 436046
rect 166048 435922 166118 435978
rect 166174 435922 166242 435978
rect 166298 435922 166368 435978
rect 166048 435888 166368 435922
rect 196768 436350 197088 436384
rect 196768 436294 196838 436350
rect 196894 436294 196962 436350
rect 197018 436294 197088 436350
rect 196768 436226 197088 436294
rect 196768 436170 196838 436226
rect 196894 436170 196962 436226
rect 197018 436170 197088 436226
rect 196768 436102 197088 436170
rect 196768 436046 196838 436102
rect 196894 436046 196962 436102
rect 197018 436046 197088 436102
rect 196768 435978 197088 436046
rect 196768 435922 196838 435978
rect 196894 435922 196962 435978
rect 197018 435922 197088 435978
rect 196768 435888 197088 435922
rect 227488 436350 227808 436384
rect 227488 436294 227558 436350
rect 227614 436294 227682 436350
rect 227738 436294 227808 436350
rect 227488 436226 227808 436294
rect 227488 436170 227558 436226
rect 227614 436170 227682 436226
rect 227738 436170 227808 436226
rect 227488 436102 227808 436170
rect 227488 436046 227558 436102
rect 227614 436046 227682 436102
rect 227738 436046 227808 436102
rect 227488 435978 227808 436046
rect 227488 435922 227558 435978
rect 227614 435922 227682 435978
rect 227738 435922 227808 435978
rect 227488 435888 227808 435922
rect 258208 436350 258528 436384
rect 258208 436294 258278 436350
rect 258334 436294 258402 436350
rect 258458 436294 258528 436350
rect 258208 436226 258528 436294
rect 258208 436170 258278 436226
rect 258334 436170 258402 436226
rect 258458 436170 258528 436226
rect 258208 436102 258528 436170
rect 258208 436046 258278 436102
rect 258334 436046 258402 436102
rect 258458 436046 258528 436102
rect 258208 435978 258528 436046
rect 258208 435922 258278 435978
rect 258334 435922 258402 435978
rect 258458 435922 258528 435978
rect 258208 435888 258528 435922
rect 288928 436350 289248 436384
rect 288928 436294 288998 436350
rect 289054 436294 289122 436350
rect 289178 436294 289248 436350
rect 288928 436226 289248 436294
rect 288928 436170 288998 436226
rect 289054 436170 289122 436226
rect 289178 436170 289248 436226
rect 288928 436102 289248 436170
rect 288928 436046 288998 436102
rect 289054 436046 289122 436102
rect 289178 436046 289248 436102
rect 288928 435978 289248 436046
rect 288928 435922 288998 435978
rect 289054 435922 289122 435978
rect 289178 435922 289248 435978
rect 288928 435888 289248 435922
rect 319648 436350 319968 436384
rect 319648 436294 319718 436350
rect 319774 436294 319842 436350
rect 319898 436294 319968 436350
rect 319648 436226 319968 436294
rect 319648 436170 319718 436226
rect 319774 436170 319842 436226
rect 319898 436170 319968 436226
rect 319648 436102 319968 436170
rect 319648 436046 319718 436102
rect 319774 436046 319842 436102
rect 319898 436046 319968 436102
rect 319648 435978 319968 436046
rect 319648 435922 319718 435978
rect 319774 435922 319842 435978
rect 319898 435922 319968 435978
rect 319648 435888 319968 435922
rect 350368 436350 350688 436384
rect 350368 436294 350438 436350
rect 350494 436294 350562 436350
rect 350618 436294 350688 436350
rect 350368 436226 350688 436294
rect 350368 436170 350438 436226
rect 350494 436170 350562 436226
rect 350618 436170 350688 436226
rect 350368 436102 350688 436170
rect 350368 436046 350438 436102
rect 350494 436046 350562 436102
rect 350618 436046 350688 436102
rect 350368 435978 350688 436046
rect 350368 435922 350438 435978
rect 350494 435922 350562 435978
rect 350618 435922 350688 435978
rect 350368 435888 350688 435922
rect 381088 436350 381408 436384
rect 381088 436294 381158 436350
rect 381214 436294 381282 436350
rect 381338 436294 381408 436350
rect 381088 436226 381408 436294
rect 381088 436170 381158 436226
rect 381214 436170 381282 436226
rect 381338 436170 381408 436226
rect 381088 436102 381408 436170
rect 381088 436046 381158 436102
rect 381214 436046 381282 436102
rect 381338 436046 381408 436102
rect 381088 435978 381408 436046
rect 381088 435922 381158 435978
rect 381214 435922 381282 435978
rect 381338 435922 381408 435978
rect 381088 435888 381408 435922
rect 411808 436350 412128 436384
rect 411808 436294 411878 436350
rect 411934 436294 412002 436350
rect 412058 436294 412128 436350
rect 411808 436226 412128 436294
rect 411808 436170 411878 436226
rect 411934 436170 412002 436226
rect 412058 436170 412128 436226
rect 411808 436102 412128 436170
rect 411808 436046 411878 436102
rect 411934 436046 412002 436102
rect 412058 436046 412128 436102
rect 411808 435978 412128 436046
rect 411808 435922 411878 435978
rect 411934 435922 412002 435978
rect 412058 435922 412128 435978
rect 411808 435888 412128 435922
rect 442528 436350 442848 436384
rect 442528 436294 442598 436350
rect 442654 436294 442722 436350
rect 442778 436294 442848 436350
rect 442528 436226 442848 436294
rect 442528 436170 442598 436226
rect 442654 436170 442722 436226
rect 442778 436170 442848 436226
rect 442528 436102 442848 436170
rect 442528 436046 442598 436102
rect 442654 436046 442722 436102
rect 442778 436046 442848 436102
rect 442528 435978 442848 436046
rect 442528 435922 442598 435978
rect 442654 435922 442722 435978
rect 442778 435922 442848 435978
rect 442528 435888 442848 435922
rect 473248 436350 473568 436384
rect 473248 436294 473318 436350
rect 473374 436294 473442 436350
rect 473498 436294 473568 436350
rect 473248 436226 473568 436294
rect 473248 436170 473318 436226
rect 473374 436170 473442 436226
rect 473498 436170 473568 436226
rect 473248 436102 473568 436170
rect 473248 436046 473318 436102
rect 473374 436046 473442 436102
rect 473498 436046 473568 436102
rect 473248 435978 473568 436046
rect 473248 435922 473318 435978
rect 473374 435922 473442 435978
rect 473498 435922 473568 435978
rect 473248 435888 473568 435922
rect 503968 436350 504288 436384
rect 503968 436294 504038 436350
rect 504094 436294 504162 436350
rect 504218 436294 504288 436350
rect 503968 436226 504288 436294
rect 503968 436170 504038 436226
rect 504094 436170 504162 436226
rect 504218 436170 504288 436226
rect 503968 436102 504288 436170
rect 503968 436046 504038 436102
rect 504094 436046 504162 436102
rect 504218 436046 504288 436102
rect 503968 435978 504288 436046
rect 503968 435922 504038 435978
rect 504094 435922 504162 435978
rect 504218 435922 504288 435978
rect 503968 435888 504288 435922
rect 534688 436350 535008 436384
rect 534688 436294 534758 436350
rect 534814 436294 534882 436350
rect 534938 436294 535008 436350
rect 534688 436226 535008 436294
rect 534688 436170 534758 436226
rect 534814 436170 534882 436226
rect 534938 436170 535008 436226
rect 534688 436102 535008 436170
rect 534688 436046 534758 436102
rect 534814 436046 534882 436102
rect 534938 436046 535008 436102
rect 534688 435978 535008 436046
rect 534688 435922 534758 435978
rect 534814 435922 534882 435978
rect 534938 435922 535008 435978
rect 534688 435888 535008 435922
rect 565408 436350 565728 436384
rect 565408 436294 565478 436350
rect 565534 436294 565602 436350
rect 565658 436294 565728 436350
rect 565408 436226 565728 436294
rect 565408 436170 565478 436226
rect 565534 436170 565602 436226
rect 565658 436170 565728 436226
rect 565408 436102 565728 436170
rect 565408 436046 565478 436102
rect 565534 436046 565602 436102
rect 565658 436046 565728 436102
rect 565408 435978 565728 436046
rect 565408 435922 565478 435978
rect 565534 435922 565602 435978
rect 565658 435922 565728 435978
rect 565408 435888 565728 435922
rect 589098 436350 589718 453922
rect 592818 460350 593438 477922
rect 592818 460294 592914 460350
rect 592970 460294 593038 460350
rect 593094 460294 593162 460350
rect 593218 460294 593286 460350
rect 593342 460294 593438 460350
rect 592818 460226 593438 460294
rect 592818 460170 592914 460226
rect 592970 460170 593038 460226
rect 593094 460170 593162 460226
rect 593218 460170 593286 460226
rect 593342 460170 593438 460226
rect 592818 460102 593438 460170
rect 592818 460046 592914 460102
rect 592970 460046 593038 460102
rect 593094 460046 593162 460102
rect 593218 460046 593286 460102
rect 593342 460046 593438 460102
rect 592818 459978 593438 460046
rect 592818 459922 592914 459978
rect 592970 459922 593038 459978
rect 593094 459922 593162 459978
rect 593218 459922 593286 459978
rect 593342 459922 593438 459978
rect 589098 436294 589194 436350
rect 589250 436294 589318 436350
rect 589374 436294 589442 436350
rect 589498 436294 589566 436350
rect 589622 436294 589718 436350
rect 589098 436226 589718 436294
rect 589098 436170 589194 436226
rect 589250 436170 589318 436226
rect 589374 436170 589442 436226
rect 589498 436170 589566 436226
rect 589622 436170 589718 436226
rect 589098 436102 589718 436170
rect 589098 436046 589194 436102
rect 589250 436046 589318 436102
rect 589374 436046 589442 436102
rect 589498 436046 589566 436102
rect 589622 436046 589718 436102
rect 589098 435978 589718 436046
rect 589098 435922 589194 435978
rect 589250 435922 589318 435978
rect 589374 435922 589442 435978
rect 589498 435922 589566 435978
rect 589622 435922 589718 435978
rect 5418 418294 5514 418350
rect 5570 418294 5638 418350
rect 5694 418294 5762 418350
rect 5818 418294 5886 418350
rect 5942 418294 6038 418350
rect 5418 418226 6038 418294
rect 5418 418170 5514 418226
rect 5570 418170 5638 418226
rect 5694 418170 5762 418226
rect 5818 418170 5886 418226
rect 5942 418170 6038 418226
rect 5418 418102 6038 418170
rect 5418 418046 5514 418102
rect 5570 418046 5638 418102
rect 5694 418046 5762 418102
rect 5818 418046 5886 418102
rect 5942 418046 6038 418102
rect 5418 417978 6038 418046
rect 5418 417922 5514 417978
rect 5570 417922 5638 417978
rect 5694 417922 5762 417978
rect 5818 417922 5886 417978
rect 5942 417922 6038 417978
rect -956 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 -336 400350
rect -956 400226 -336 400294
rect -956 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 -336 400226
rect -956 400102 -336 400170
rect -956 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 -336 400102
rect -956 399978 -336 400046
rect -956 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 -336 399978
rect -956 382350 -336 399922
rect 4172 403732 4228 403742
rect 4172 386148 4228 403676
rect 4172 386082 4228 386092
rect 5418 400350 6038 417922
rect 6412 431956 6468 431966
rect 5418 400294 5514 400350
rect 5570 400294 5638 400350
rect 5694 400294 5762 400350
rect 5818 400294 5886 400350
rect 5942 400294 6038 400350
rect 5418 400226 6038 400294
rect 5418 400170 5514 400226
rect 5570 400170 5638 400226
rect 5694 400170 5762 400226
rect 5818 400170 5886 400226
rect 5942 400170 6038 400226
rect 5418 400102 6038 400170
rect 5418 400046 5514 400102
rect 5570 400046 5638 400102
rect 5694 400046 5762 400102
rect 5818 400046 5886 400102
rect 5942 400046 6038 400102
rect 5418 399978 6038 400046
rect 5418 399922 5514 399978
rect 5570 399922 5638 399978
rect 5694 399922 5762 399978
rect 5818 399922 5886 399978
rect 5942 399922 6038 399978
rect -956 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 -336 382350
rect -956 382226 -336 382294
rect -956 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 -336 382226
rect -956 382102 -336 382170
rect -956 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 -336 382102
rect -956 381978 -336 382046
rect -956 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 -336 381978
rect -956 364350 -336 381922
rect -956 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 -336 364350
rect -956 364226 -336 364294
rect -956 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 -336 364226
rect -956 364102 -336 364170
rect -956 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 -336 364102
rect -956 363978 -336 364046
rect -956 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 -336 363978
rect -956 346350 -336 363922
rect 5418 382350 6038 399922
rect 6188 417844 6244 417854
rect 6188 396676 6244 417788
rect 6412 417732 6468 431900
rect 585452 430164 585508 430174
rect 27808 424350 28128 424384
rect 27808 424294 27878 424350
rect 27934 424294 28002 424350
rect 28058 424294 28128 424350
rect 27808 424226 28128 424294
rect 27808 424170 27878 424226
rect 27934 424170 28002 424226
rect 28058 424170 28128 424226
rect 27808 424102 28128 424170
rect 27808 424046 27878 424102
rect 27934 424046 28002 424102
rect 28058 424046 28128 424102
rect 27808 423978 28128 424046
rect 27808 423922 27878 423978
rect 27934 423922 28002 423978
rect 28058 423922 28128 423978
rect 27808 423888 28128 423922
rect 58528 424350 58848 424384
rect 58528 424294 58598 424350
rect 58654 424294 58722 424350
rect 58778 424294 58848 424350
rect 58528 424226 58848 424294
rect 58528 424170 58598 424226
rect 58654 424170 58722 424226
rect 58778 424170 58848 424226
rect 58528 424102 58848 424170
rect 58528 424046 58598 424102
rect 58654 424046 58722 424102
rect 58778 424046 58848 424102
rect 58528 423978 58848 424046
rect 58528 423922 58598 423978
rect 58654 423922 58722 423978
rect 58778 423922 58848 423978
rect 58528 423888 58848 423922
rect 89248 424350 89568 424384
rect 89248 424294 89318 424350
rect 89374 424294 89442 424350
rect 89498 424294 89568 424350
rect 89248 424226 89568 424294
rect 89248 424170 89318 424226
rect 89374 424170 89442 424226
rect 89498 424170 89568 424226
rect 89248 424102 89568 424170
rect 89248 424046 89318 424102
rect 89374 424046 89442 424102
rect 89498 424046 89568 424102
rect 89248 423978 89568 424046
rect 89248 423922 89318 423978
rect 89374 423922 89442 423978
rect 89498 423922 89568 423978
rect 89248 423888 89568 423922
rect 119968 424350 120288 424384
rect 119968 424294 120038 424350
rect 120094 424294 120162 424350
rect 120218 424294 120288 424350
rect 119968 424226 120288 424294
rect 119968 424170 120038 424226
rect 120094 424170 120162 424226
rect 120218 424170 120288 424226
rect 119968 424102 120288 424170
rect 119968 424046 120038 424102
rect 120094 424046 120162 424102
rect 120218 424046 120288 424102
rect 119968 423978 120288 424046
rect 119968 423922 120038 423978
rect 120094 423922 120162 423978
rect 120218 423922 120288 423978
rect 119968 423888 120288 423922
rect 150688 424350 151008 424384
rect 150688 424294 150758 424350
rect 150814 424294 150882 424350
rect 150938 424294 151008 424350
rect 150688 424226 151008 424294
rect 150688 424170 150758 424226
rect 150814 424170 150882 424226
rect 150938 424170 151008 424226
rect 150688 424102 151008 424170
rect 150688 424046 150758 424102
rect 150814 424046 150882 424102
rect 150938 424046 151008 424102
rect 150688 423978 151008 424046
rect 150688 423922 150758 423978
rect 150814 423922 150882 423978
rect 150938 423922 151008 423978
rect 150688 423888 151008 423922
rect 181408 424350 181728 424384
rect 181408 424294 181478 424350
rect 181534 424294 181602 424350
rect 181658 424294 181728 424350
rect 181408 424226 181728 424294
rect 181408 424170 181478 424226
rect 181534 424170 181602 424226
rect 181658 424170 181728 424226
rect 181408 424102 181728 424170
rect 181408 424046 181478 424102
rect 181534 424046 181602 424102
rect 181658 424046 181728 424102
rect 181408 423978 181728 424046
rect 181408 423922 181478 423978
rect 181534 423922 181602 423978
rect 181658 423922 181728 423978
rect 181408 423888 181728 423922
rect 212128 424350 212448 424384
rect 212128 424294 212198 424350
rect 212254 424294 212322 424350
rect 212378 424294 212448 424350
rect 212128 424226 212448 424294
rect 212128 424170 212198 424226
rect 212254 424170 212322 424226
rect 212378 424170 212448 424226
rect 212128 424102 212448 424170
rect 212128 424046 212198 424102
rect 212254 424046 212322 424102
rect 212378 424046 212448 424102
rect 212128 423978 212448 424046
rect 212128 423922 212198 423978
rect 212254 423922 212322 423978
rect 212378 423922 212448 423978
rect 212128 423888 212448 423922
rect 242848 424350 243168 424384
rect 242848 424294 242918 424350
rect 242974 424294 243042 424350
rect 243098 424294 243168 424350
rect 242848 424226 243168 424294
rect 242848 424170 242918 424226
rect 242974 424170 243042 424226
rect 243098 424170 243168 424226
rect 242848 424102 243168 424170
rect 242848 424046 242918 424102
rect 242974 424046 243042 424102
rect 243098 424046 243168 424102
rect 242848 423978 243168 424046
rect 242848 423922 242918 423978
rect 242974 423922 243042 423978
rect 243098 423922 243168 423978
rect 242848 423888 243168 423922
rect 273568 424350 273888 424384
rect 273568 424294 273638 424350
rect 273694 424294 273762 424350
rect 273818 424294 273888 424350
rect 273568 424226 273888 424294
rect 273568 424170 273638 424226
rect 273694 424170 273762 424226
rect 273818 424170 273888 424226
rect 273568 424102 273888 424170
rect 273568 424046 273638 424102
rect 273694 424046 273762 424102
rect 273818 424046 273888 424102
rect 273568 423978 273888 424046
rect 273568 423922 273638 423978
rect 273694 423922 273762 423978
rect 273818 423922 273888 423978
rect 273568 423888 273888 423922
rect 304288 424350 304608 424384
rect 304288 424294 304358 424350
rect 304414 424294 304482 424350
rect 304538 424294 304608 424350
rect 304288 424226 304608 424294
rect 304288 424170 304358 424226
rect 304414 424170 304482 424226
rect 304538 424170 304608 424226
rect 304288 424102 304608 424170
rect 304288 424046 304358 424102
rect 304414 424046 304482 424102
rect 304538 424046 304608 424102
rect 304288 423978 304608 424046
rect 304288 423922 304358 423978
rect 304414 423922 304482 423978
rect 304538 423922 304608 423978
rect 304288 423888 304608 423922
rect 335008 424350 335328 424384
rect 335008 424294 335078 424350
rect 335134 424294 335202 424350
rect 335258 424294 335328 424350
rect 335008 424226 335328 424294
rect 335008 424170 335078 424226
rect 335134 424170 335202 424226
rect 335258 424170 335328 424226
rect 335008 424102 335328 424170
rect 335008 424046 335078 424102
rect 335134 424046 335202 424102
rect 335258 424046 335328 424102
rect 335008 423978 335328 424046
rect 335008 423922 335078 423978
rect 335134 423922 335202 423978
rect 335258 423922 335328 423978
rect 335008 423888 335328 423922
rect 365728 424350 366048 424384
rect 365728 424294 365798 424350
rect 365854 424294 365922 424350
rect 365978 424294 366048 424350
rect 365728 424226 366048 424294
rect 365728 424170 365798 424226
rect 365854 424170 365922 424226
rect 365978 424170 366048 424226
rect 365728 424102 366048 424170
rect 365728 424046 365798 424102
rect 365854 424046 365922 424102
rect 365978 424046 366048 424102
rect 365728 423978 366048 424046
rect 365728 423922 365798 423978
rect 365854 423922 365922 423978
rect 365978 423922 366048 423978
rect 365728 423888 366048 423922
rect 396448 424350 396768 424384
rect 396448 424294 396518 424350
rect 396574 424294 396642 424350
rect 396698 424294 396768 424350
rect 396448 424226 396768 424294
rect 396448 424170 396518 424226
rect 396574 424170 396642 424226
rect 396698 424170 396768 424226
rect 396448 424102 396768 424170
rect 396448 424046 396518 424102
rect 396574 424046 396642 424102
rect 396698 424046 396768 424102
rect 396448 423978 396768 424046
rect 396448 423922 396518 423978
rect 396574 423922 396642 423978
rect 396698 423922 396768 423978
rect 396448 423888 396768 423922
rect 427168 424350 427488 424384
rect 427168 424294 427238 424350
rect 427294 424294 427362 424350
rect 427418 424294 427488 424350
rect 427168 424226 427488 424294
rect 427168 424170 427238 424226
rect 427294 424170 427362 424226
rect 427418 424170 427488 424226
rect 427168 424102 427488 424170
rect 427168 424046 427238 424102
rect 427294 424046 427362 424102
rect 427418 424046 427488 424102
rect 427168 423978 427488 424046
rect 427168 423922 427238 423978
rect 427294 423922 427362 423978
rect 427418 423922 427488 423978
rect 427168 423888 427488 423922
rect 457888 424350 458208 424384
rect 457888 424294 457958 424350
rect 458014 424294 458082 424350
rect 458138 424294 458208 424350
rect 457888 424226 458208 424294
rect 457888 424170 457958 424226
rect 458014 424170 458082 424226
rect 458138 424170 458208 424226
rect 457888 424102 458208 424170
rect 457888 424046 457958 424102
rect 458014 424046 458082 424102
rect 458138 424046 458208 424102
rect 457888 423978 458208 424046
rect 457888 423922 457958 423978
rect 458014 423922 458082 423978
rect 458138 423922 458208 423978
rect 457888 423888 458208 423922
rect 488608 424350 488928 424384
rect 488608 424294 488678 424350
rect 488734 424294 488802 424350
rect 488858 424294 488928 424350
rect 488608 424226 488928 424294
rect 488608 424170 488678 424226
rect 488734 424170 488802 424226
rect 488858 424170 488928 424226
rect 488608 424102 488928 424170
rect 488608 424046 488678 424102
rect 488734 424046 488802 424102
rect 488858 424046 488928 424102
rect 488608 423978 488928 424046
rect 488608 423922 488678 423978
rect 488734 423922 488802 423978
rect 488858 423922 488928 423978
rect 488608 423888 488928 423922
rect 519328 424350 519648 424384
rect 519328 424294 519398 424350
rect 519454 424294 519522 424350
rect 519578 424294 519648 424350
rect 519328 424226 519648 424294
rect 519328 424170 519398 424226
rect 519454 424170 519522 424226
rect 519578 424170 519648 424226
rect 519328 424102 519648 424170
rect 519328 424046 519398 424102
rect 519454 424046 519522 424102
rect 519578 424046 519648 424102
rect 519328 423978 519648 424046
rect 519328 423922 519398 423978
rect 519454 423922 519522 423978
rect 519578 423922 519648 423978
rect 519328 423888 519648 423922
rect 550048 424350 550368 424384
rect 550048 424294 550118 424350
rect 550174 424294 550242 424350
rect 550298 424294 550368 424350
rect 550048 424226 550368 424294
rect 550048 424170 550118 424226
rect 550174 424170 550242 424226
rect 550298 424170 550368 424226
rect 550048 424102 550368 424170
rect 550048 424046 550118 424102
rect 550174 424046 550242 424102
rect 550298 424046 550368 424102
rect 550048 423978 550368 424046
rect 550048 423922 550118 423978
rect 550174 423922 550242 423978
rect 550298 423922 550368 423978
rect 550048 423888 550368 423922
rect 12448 418350 12768 418384
rect 12448 418294 12518 418350
rect 12574 418294 12642 418350
rect 12698 418294 12768 418350
rect 12448 418226 12768 418294
rect 12448 418170 12518 418226
rect 12574 418170 12642 418226
rect 12698 418170 12768 418226
rect 12448 418102 12768 418170
rect 12448 418046 12518 418102
rect 12574 418046 12642 418102
rect 12698 418046 12768 418102
rect 12448 417978 12768 418046
rect 12448 417922 12518 417978
rect 12574 417922 12642 417978
rect 12698 417922 12768 417978
rect 12448 417888 12768 417922
rect 43168 418350 43488 418384
rect 43168 418294 43238 418350
rect 43294 418294 43362 418350
rect 43418 418294 43488 418350
rect 43168 418226 43488 418294
rect 43168 418170 43238 418226
rect 43294 418170 43362 418226
rect 43418 418170 43488 418226
rect 43168 418102 43488 418170
rect 43168 418046 43238 418102
rect 43294 418046 43362 418102
rect 43418 418046 43488 418102
rect 43168 417978 43488 418046
rect 43168 417922 43238 417978
rect 43294 417922 43362 417978
rect 43418 417922 43488 417978
rect 43168 417888 43488 417922
rect 73888 418350 74208 418384
rect 73888 418294 73958 418350
rect 74014 418294 74082 418350
rect 74138 418294 74208 418350
rect 73888 418226 74208 418294
rect 73888 418170 73958 418226
rect 74014 418170 74082 418226
rect 74138 418170 74208 418226
rect 73888 418102 74208 418170
rect 73888 418046 73958 418102
rect 74014 418046 74082 418102
rect 74138 418046 74208 418102
rect 73888 417978 74208 418046
rect 73888 417922 73958 417978
rect 74014 417922 74082 417978
rect 74138 417922 74208 417978
rect 73888 417888 74208 417922
rect 104608 418350 104928 418384
rect 104608 418294 104678 418350
rect 104734 418294 104802 418350
rect 104858 418294 104928 418350
rect 104608 418226 104928 418294
rect 104608 418170 104678 418226
rect 104734 418170 104802 418226
rect 104858 418170 104928 418226
rect 104608 418102 104928 418170
rect 104608 418046 104678 418102
rect 104734 418046 104802 418102
rect 104858 418046 104928 418102
rect 104608 417978 104928 418046
rect 104608 417922 104678 417978
rect 104734 417922 104802 417978
rect 104858 417922 104928 417978
rect 104608 417888 104928 417922
rect 135328 418350 135648 418384
rect 135328 418294 135398 418350
rect 135454 418294 135522 418350
rect 135578 418294 135648 418350
rect 135328 418226 135648 418294
rect 135328 418170 135398 418226
rect 135454 418170 135522 418226
rect 135578 418170 135648 418226
rect 135328 418102 135648 418170
rect 135328 418046 135398 418102
rect 135454 418046 135522 418102
rect 135578 418046 135648 418102
rect 135328 417978 135648 418046
rect 135328 417922 135398 417978
rect 135454 417922 135522 417978
rect 135578 417922 135648 417978
rect 135328 417888 135648 417922
rect 166048 418350 166368 418384
rect 166048 418294 166118 418350
rect 166174 418294 166242 418350
rect 166298 418294 166368 418350
rect 166048 418226 166368 418294
rect 166048 418170 166118 418226
rect 166174 418170 166242 418226
rect 166298 418170 166368 418226
rect 166048 418102 166368 418170
rect 166048 418046 166118 418102
rect 166174 418046 166242 418102
rect 166298 418046 166368 418102
rect 166048 417978 166368 418046
rect 166048 417922 166118 417978
rect 166174 417922 166242 417978
rect 166298 417922 166368 417978
rect 166048 417888 166368 417922
rect 196768 418350 197088 418384
rect 196768 418294 196838 418350
rect 196894 418294 196962 418350
rect 197018 418294 197088 418350
rect 196768 418226 197088 418294
rect 196768 418170 196838 418226
rect 196894 418170 196962 418226
rect 197018 418170 197088 418226
rect 196768 418102 197088 418170
rect 196768 418046 196838 418102
rect 196894 418046 196962 418102
rect 197018 418046 197088 418102
rect 196768 417978 197088 418046
rect 196768 417922 196838 417978
rect 196894 417922 196962 417978
rect 197018 417922 197088 417978
rect 196768 417888 197088 417922
rect 227488 418350 227808 418384
rect 227488 418294 227558 418350
rect 227614 418294 227682 418350
rect 227738 418294 227808 418350
rect 227488 418226 227808 418294
rect 227488 418170 227558 418226
rect 227614 418170 227682 418226
rect 227738 418170 227808 418226
rect 227488 418102 227808 418170
rect 227488 418046 227558 418102
rect 227614 418046 227682 418102
rect 227738 418046 227808 418102
rect 227488 417978 227808 418046
rect 227488 417922 227558 417978
rect 227614 417922 227682 417978
rect 227738 417922 227808 417978
rect 227488 417888 227808 417922
rect 258208 418350 258528 418384
rect 258208 418294 258278 418350
rect 258334 418294 258402 418350
rect 258458 418294 258528 418350
rect 258208 418226 258528 418294
rect 258208 418170 258278 418226
rect 258334 418170 258402 418226
rect 258458 418170 258528 418226
rect 258208 418102 258528 418170
rect 258208 418046 258278 418102
rect 258334 418046 258402 418102
rect 258458 418046 258528 418102
rect 258208 417978 258528 418046
rect 258208 417922 258278 417978
rect 258334 417922 258402 417978
rect 258458 417922 258528 417978
rect 258208 417888 258528 417922
rect 288928 418350 289248 418384
rect 288928 418294 288998 418350
rect 289054 418294 289122 418350
rect 289178 418294 289248 418350
rect 288928 418226 289248 418294
rect 288928 418170 288998 418226
rect 289054 418170 289122 418226
rect 289178 418170 289248 418226
rect 288928 418102 289248 418170
rect 288928 418046 288998 418102
rect 289054 418046 289122 418102
rect 289178 418046 289248 418102
rect 288928 417978 289248 418046
rect 288928 417922 288998 417978
rect 289054 417922 289122 417978
rect 289178 417922 289248 417978
rect 288928 417888 289248 417922
rect 319648 418350 319968 418384
rect 319648 418294 319718 418350
rect 319774 418294 319842 418350
rect 319898 418294 319968 418350
rect 319648 418226 319968 418294
rect 319648 418170 319718 418226
rect 319774 418170 319842 418226
rect 319898 418170 319968 418226
rect 319648 418102 319968 418170
rect 319648 418046 319718 418102
rect 319774 418046 319842 418102
rect 319898 418046 319968 418102
rect 319648 417978 319968 418046
rect 319648 417922 319718 417978
rect 319774 417922 319842 417978
rect 319898 417922 319968 417978
rect 319648 417888 319968 417922
rect 350368 418350 350688 418384
rect 350368 418294 350438 418350
rect 350494 418294 350562 418350
rect 350618 418294 350688 418350
rect 350368 418226 350688 418294
rect 350368 418170 350438 418226
rect 350494 418170 350562 418226
rect 350618 418170 350688 418226
rect 350368 418102 350688 418170
rect 350368 418046 350438 418102
rect 350494 418046 350562 418102
rect 350618 418046 350688 418102
rect 350368 417978 350688 418046
rect 350368 417922 350438 417978
rect 350494 417922 350562 417978
rect 350618 417922 350688 417978
rect 350368 417888 350688 417922
rect 381088 418350 381408 418384
rect 381088 418294 381158 418350
rect 381214 418294 381282 418350
rect 381338 418294 381408 418350
rect 381088 418226 381408 418294
rect 381088 418170 381158 418226
rect 381214 418170 381282 418226
rect 381338 418170 381408 418226
rect 381088 418102 381408 418170
rect 381088 418046 381158 418102
rect 381214 418046 381282 418102
rect 381338 418046 381408 418102
rect 381088 417978 381408 418046
rect 381088 417922 381158 417978
rect 381214 417922 381282 417978
rect 381338 417922 381408 417978
rect 381088 417888 381408 417922
rect 411808 418350 412128 418384
rect 411808 418294 411878 418350
rect 411934 418294 412002 418350
rect 412058 418294 412128 418350
rect 411808 418226 412128 418294
rect 411808 418170 411878 418226
rect 411934 418170 412002 418226
rect 412058 418170 412128 418226
rect 411808 418102 412128 418170
rect 411808 418046 411878 418102
rect 411934 418046 412002 418102
rect 412058 418046 412128 418102
rect 411808 417978 412128 418046
rect 411808 417922 411878 417978
rect 411934 417922 412002 417978
rect 412058 417922 412128 417978
rect 411808 417888 412128 417922
rect 442528 418350 442848 418384
rect 442528 418294 442598 418350
rect 442654 418294 442722 418350
rect 442778 418294 442848 418350
rect 442528 418226 442848 418294
rect 442528 418170 442598 418226
rect 442654 418170 442722 418226
rect 442778 418170 442848 418226
rect 442528 418102 442848 418170
rect 442528 418046 442598 418102
rect 442654 418046 442722 418102
rect 442778 418046 442848 418102
rect 442528 417978 442848 418046
rect 442528 417922 442598 417978
rect 442654 417922 442722 417978
rect 442778 417922 442848 417978
rect 442528 417888 442848 417922
rect 473248 418350 473568 418384
rect 473248 418294 473318 418350
rect 473374 418294 473442 418350
rect 473498 418294 473568 418350
rect 473248 418226 473568 418294
rect 473248 418170 473318 418226
rect 473374 418170 473442 418226
rect 473498 418170 473568 418226
rect 473248 418102 473568 418170
rect 473248 418046 473318 418102
rect 473374 418046 473442 418102
rect 473498 418046 473568 418102
rect 473248 417978 473568 418046
rect 473248 417922 473318 417978
rect 473374 417922 473442 417978
rect 473498 417922 473568 417978
rect 473248 417888 473568 417922
rect 503968 418350 504288 418384
rect 503968 418294 504038 418350
rect 504094 418294 504162 418350
rect 504218 418294 504288 418350
rect 503968 418226 504288 418294
rect 503968 418170 504038 418226
rect 504094 418170 504162 418226
rect 504218 418170 504288 418226
rect 503968 418102 504288 418170
rect 503968 418046 504038 418102
rect 504094 418046 504162 418102
rect 504218 418046 504288 418102
rect 503968 417978 504288 418046
rect 503968 417922 504038 417978
rect 504094 417922 504162 417978
rect 504218 417922 504288 417978
rect 503968 417888 504288 417922
rect 534688 418350 535008 418384
rect 534688 418294 534758 418350
rect 534814 418294 534882 418350
rect 534938 418294 535008 418350
rect 534688 418226 535008 418294
rect 534688 418170 534758 418226
rect 534814 418170 534882 418226
rect 534938 418170 535008 418226
rect 534688 418102 535008 418170
rect 534688 418046 534758 418102
rect 534814 418046 534882 418102
rect 534938 418046 535008 418102
rect 534688 417978 535008 418046
rect 534688 417922 534758 417978
rect 534814 417922 534882 417978
rect 534938 417922 535008 417978
rect 534688 417888 535008 417922
rect 565408 418350 565728 418384
rect 565408 418294 565478 418350
rect 565534 418294 565602 418350
rect 565658 418294 565728 418350
rect 565408 418226 565728 418294
rect 565408 418170 565478 418226
rect 565534 418170 565602 418226
rect 565658 418170 565728 418226
rect 565408 418102 565728 418170
rect 565408 418046 565478 418102
rect 565534 418046 565602 418102
rect 565658 418046 565728 418102
rect 565408 417978 565728 418046
rect 565408 417922 565478 417978
rect 565534 417922 565602 417978
rect 565658 417922 565728 417978
rect 565408 417888 565728 417922
rect 6412 417666 6468 417676
rect 27808 406350 28128 406384
rect 27808 406294 27878 406350
rect 27934 406294 28002 406350
rect 28058 406294 28128 406350
rect 27808 406226 28128 406294
rect 27808 406170 27878 406226
rect 27934 406170 28002 406226
rect 28058 406170 28128 406226
rect 27808 406102 28128 406170
rect 27808 406046 27878 406102
rect 27934 406046 28002 406102
rect 28058 406046 28128 406102
rect 27808 405978 28128 406046
rect 27808 405922 27878 405978
rect 27934 405922 28002 405978
rect 28058 405922 28128 405978
rect 27808 405888 28128 405922
rect 58528 406350 58848 406384
rect 58528 406294 58598 406350
rect 58654 406294 58722 406350
rect 58778 406294 58848 406350
rect 58528 406226 58848 406294
rect 58528 406170 58598 406226
rect 58654 406170 58722 406226
rect 58778 406170 58848 406226
rect 58528 406102 58848 406170
rect 58528 406046 58598 406102
rect 58654 406046 58722 406102
rect 58778 406046 58848 406102
rect 58528 405978 58848 406046
rect 58528 405922 58598 405978
rect 58654 405922 58722 405978
rect 58778 405922 58848 405978
rect 58528 405888 58848 405922
rect 89248 406350 89568 406384
rect 89248 406294 89318 406350
rect 89374 406294 89442 406350
rect 89498 406294 89568 406350
rect 89248 406226 89568 406294
rect 89248 406170 89318 406226
rect 89374 406170 89442 406226
rect 89498 406170 89568 406226
rect 89248 406102 89568 406170
rect 89248 406046 89318 406102
rect 89374 406046 89442 406102
rect 89498 406046 89568 406102
rect 89248 405978 89568 406046
rect 89248 405922 89318 405978
rect 89374 405922 89442 405978
rect 89498 405922 89568 405978
rect 89248 405888 89568 405922
rect 119968 406350 120288 406384
rect 119968 406294 120038 406350
rect 120094 406294 120162 406350
rect 120218 406294 120288 406350
rect 119968 406226 120288 406294
rect 119968 406170 120038 406226
rect 120094 406170 120162 406226
rect 120218 406170 120288 406226
rect 119968 406102 120288 406170
rect 119968 406046 120038 406102
rect 120094 406046 120162 406102
rect 120218 406046 120288 406102
rect 119968 405978 120288 406046
rect 119968 405922 120038 405978
rect 120094 405922 120162 405978
rect 120218 405922 120288 405978
rect 119968 405888 120288 405922
rect 150688 406350 151008 406384
rect 150688 406294 150758 406350
rect 150814 406294 150882 406350
rect 150938 406294 151008 406350
rect 150688 406226 151008 406294
rect 150688 406170 150758 406226
rect 150814 406170 150882 406226
rect 150938 406170 151008 406226
rect 150688 406102 151008 406170
rect 150688 406046 150758 406102
rect 150814 406046 150882 406102
rect 150938 406046 151008 406102
rect 150688 405978 151008 406046
rect 150688 405922 150758 405978
rect 150814 405922 150882 405978
rect 150938 405922 151008 405978
rect 150688 405888 151008 405922
rect 181408 406350 181728 406384
rect 181408 406294 181478 406350
rect 181534 406294 181602 406350
rect 181658 406294 181728 406350
rect 181408 406226 181728 406294
rect 181408 406170 181478 406226
rect 181534 406170 181602 406226
rect 181658 406170 181728 406226
rect 181408 406102 181728 406170
rect 181408 406046 181478 406102
rect 181534 406046 181602 406102
rect 181658 406046 181728 406102
rect 181408 405978 181728 406046
rect 181408 405922 181478 405978
rect 181534 405922 181602 405978
rect 181658 405922 181728 405978
rect 181408 405888 181728 405922
rect 212128 406350 212448 406384
rect 212128 406294 212198 406350
rect 212254 406294 212322 406350
rect 212378 406294 212448 406350
rect 212128 406226 212448 406294
rect 212128 406170 212198 406226
rect 212254 406170 212322 406226
rect 212378 406170 212448 406226
rect 212128 406102 212448 406170
rect 212128 406046 212198 406102
rect 212254 406046 212322 406102
rect 212378 406046 212448 406102
rect 212128 405978 212448 406046
rect 212128 405922 212198 405978
rect 212254 405922 212322 405978
rect 212378 405922 212448 405978
rect 212128 405888 212448 405922
rect 242848 406350 243168 406384
rect 242848 406294 242918 406350
rect 242974 406294 243042 406350
rect 243098 406294 243168 406350
rect 242848 406226 243168 406294
rect 242848 406170 242918 406226
rect 242974 406170 243042 406226
rect 243098 406170 243168 406226
rect 242848 406102 243168 406170
rect 242848 406046 242918 406102
rect 242974 406046 243042 406102
rect 243098 406046 243168 406102
rect 242848 405978 243168 406046
rect 242848 405922 242918 405978
rect 242974 405922 243042 405978
rect 243098 405922 243168 405978
rect 242848 405888 243168 405922
rect 273568 406350 273888 406384
rect 273568 406294 273638 406350
rect 273694 406294 273762 406350
rect 273818 406294 273888 406350
rect 273568 406226 273888 406294
rect 273568 406170 273638 406226
rect 273694 406170 273762 406226
rect 273818 406170 273888 406226
rect 273568 406102 273888 406170
rect 273568 406046 273638 406102
rect 273694 406046 273762 406102
rect 273818 406046 273888 406102
rect 273568 405978 273888 406046
rect 273568 405922 273638 405978
rect 273694 405922 273762 405978
rect 273818 405922 273888 405978
rect 273568 405888 273888 405922
rect 304288 406350 304608 406384
rect 304288 406294 304358 406350
rect 304414 406294 304482 406350
rect 304538 406294 304608 406350
rect 304288 406226 304608 406294
rect 304288 406170 304358 406226
rect 304414 406170 304482 406226
rect 304538 406170 304608 406226
rect 304288 406102 304608 406170
rect 304288 406046 304358 406102
rect 304414 406046 304482 406102
rect 304538 406046 304608 406102
rect 304288 405978 304608 406046
rect 304288 405922 304358 405978
rect 304414 405922 304482 405978
rect 304538 405922 304608 405978
rect 304288 405888 304608 405922
rect 335008 406350 335328 406384
rect 335008 406294 335078 406350
rect 335134 406294 335202 406350
rect 335258 406294 335328 406350
rect 335008 406226 335328 406294
rect 335008 406170 335078 406226
rect 335134 406170 335202 406226
rect 335258 406170 335328 406226
rect 335008 406102 335328 406170
rect 335008 406046 335078 406102
rect 335134 406046 335202 406102
rect 335258 406046 335328 406102
rect 335008 405978 335328 406046
rect 335008 405922 335078 405978
rect 335134 405922 335202 405978
rect 335258 405922 335328 405978
rect 335008 405888 335328 405922
rect 365728 406350 366048 406384
rect 365728 406294 365798 406350
rect 365854 406294 365922 406350
rect 365978 406294 366048 406350
rect 365728 406226 366048 406294
rect 365728 406170 365798 406226
rect 365854 406170 365922 406226
rect 365978 406170 366048 406226
rect 365728 406102 366048 406170
rect 365728 406046 365798 406102
rect 365854 406046 365922 406102
rect 365978 406046 366048 406102
rect 365728 405978 366048 406046
rect 365728 405922 365798 405978
rect 365854 405922 365922 405978
rect 365978 405922 366048 405978
rect 365728 405888 366048 405922
rect 396448 406350 396768 406384
rect 396448 406294 396518 406350
rect 396574 406294 396642 406350
rect 396698 406294 396768 406350
rect 396448 406226 396768 406294
rect 396448 406170 396518 406226
rect 396574 406170 396642 406226
rect 396698 406170 396768 406226
rect 396448 406102 396768 406170
rect 396448 406046 396518 406102
rect 396574 406046 396642 406102
rect 396698 406046 396768 406102
rect 396448 405978 396768 406046
rect 396448 405922 396518 405978
rect 396574 405922 396642 405978
rect 396698 405922 396768 405978
rect 396448 405888 396768 405922
rect 427168 406350 427488 406384
rect 427168 406294 427238 406350
rect 427294 406294 427362 406350
rect 427418 406294 427488 406350
rect 427168 406226 427488 406294
rect 427168 406170 427238 406226
rect 427294 406170 427362 406226
rect 427418 406170 427488 406226
rect 427168 406102 427488 406170
rect 427168 406046 427238 406102
rect 427294 406046 427362 406102
rect 427418 406046 427488 406102
rect 427168 405978 427488 406046
rect 427168 405922 427238 405978
rect 427294 405922 427362 405978
rect 427418 405922 427488 405978
rect 427168 405888 427488 405922
rect 457888 406350 458208 406384
rect 457888 406294 457958 406350
rect 458014 406294 458082 406350
rect 458138 406294 458208 406350
rect 457888 406226 458208 406294
rect 457888 406170 457958 406226
rect 458014 406170 458082 406226
rect 458138 406170 458208 406226
rect 457888 406102 458208 406170
rect 457888 406046 457958 406102
rect 458014 406046 458082 406102
rect 458138 406046 458208 406102
rect 457888 405978 458208 406046
rect 457888 405922 457958 405978
rect 458014 405922 458082 405978
rect 458138 405922 458208 405978
rect 457888 405888 458208 405922
rect 488608 406350 488928 406384
rect 488608 406294 488678 406350
rect 488734 406294 488802 406350
rect 488858 406294 488928 406350
rect 488608 406226 488928 406294
rect 488608 406170 488678 406226
rect 488734 406170 488802 406226
rect 488858 406170 488928 406226
rect 488608 406102 488928 406170
rect 488608 406046 488678 406102
rect 488734 406046 488802 406102
rect 488858 406046 488928 406102
rect 488608 405978 488928 406046
rect 488608 405922 488678 405978
rect 488734 405922 488802 405978
rect 488858 405922 488928 405978
rect 488608 405888 488928 405922
rect 519328 406350 519648 406384
rect 519328 406294 519398 406350
rect 519454 406294 519522 406350
rect 519578 406294 519648 406350
rect 519328 406226 519648 406294
rect 519328 406170 519398 406226
rect 519454 406170 519522 406226
rect 519578 406170 519648 406226
rect 519328 406102 519648 406170
rect 519328 406046 519398 406102
rect 519454 406046 519522 406102
rect 519578 406046 519648 406102
rect 519328 405978 519648 406046
rect 519328 405922 519398 405978
rect 519454 405922 519522 405978
rect 519578 405922 519648 405978
rect 519328 405888 519648 405922
rect 550048 406350 550368 406384
rect 550048 406294 550118 406350
rect 550174 406294 550242 406350
rect 550298 406294 550368 406350
rect 550048 406226 550368 406294
rect 550048 406170 550118 406226
rect 550174 406170 550242 406226
rect 550298 406170 550368 406226
rect 550048 406102 550368 406170
rect 550048 406046 550118 406102
rect 550174 406046 550242 406102
rect 550298 406046 550368 406102
rect 550048 405978 550368 406046
rect 550048 405922 550118 405978
rect 550174 405922 550242 405978
rect 550298 405922 550368 405978
rect 550048 405888 550368 405922
rect 585452 404292 585508 430108
rect 589098 418350 589718 435922
rect 590492 443268 590548 443278
rect 590492 425796 590548 443212
rect 590492 425730 590548 425740
rect 592818 442350 593438 459922
rect 592818 442294 592914 442350
rect 592970 442294 593038 442350
rect 593094 442294 593162 442350
rect 593218 442294 593286 442350
rect 593342 442294 593438 442350
rect 592818 442226 593438 442294
rect 592818 442170 592914 442226
rect 592970 442170 593038 442226
rect 593094 442170 593162 442226
rect 593218 442170 593286 442226
rect 593342 442170 593438 442226
rect 592818 442102 593438 442170
rect 592818 442046 592914 442102
rect 592970 442046 593038 442102
rect 593094 442046 593162 442102
rect 593218 442046 593286 442102
rect 593342 442046 593438 442102
rect 592818 441978 593438 442046
rect 592818 441922 592914 441978
rect 592970 441922 593038 441978
rect 593094 441922 593162 441978
rect 593218 441922 593286 441978
rect 593342 441922 593438 441978
rect 589098 418294 589194 418350
rect 589250 418294 589318 418350
rect 589374 418294 589442 418350
rect 589498 418294 589566 418350
rect 589622 418294 589718 418350
rect 589098 418226 589718 418294
rect 589098 418170 589194 418226
rect 589250 418170 589318 418226
rect 589374 418170 589442 418226
rect 589498 418170 589566 418226
rect 589622 418170 589718 418226
rect 589098 418102 589718 418170
rect 589098 418046 589194 418102
rect 589250 418046 589318 418102
rect 589374 418046 589442 418102
rect 589498 418046 589566 418102
rect 589622 418046 589718 418102
rect 589098 417978 589718 418046
rect 589098 417922 589194 417978
rect 589250 417922 589318 417978
rect 589374 417922 589442 417978
rect 589498 417922 589566 417978
rect 589622 417922 589718 417978
rect 585452 404226 585508 404236
rect 585564 416836 585620 416846
rect 12448 400350 12768 400384
rect 12448 400294 12518 400350
rect 12574 400294 12642 400350
rect 12698 400294 12768 400350
rect 12448 400226 12768 400294
rect 12448 400170 12518 400226
rect 12574 400170 12642 400226
rect 12698 400170 12768 400226
rect 12448 400102 12768 400170
rect 12448 400046 12518 400102
rect 12574 400046 12642 400102
rect 12698 400046 12768 400102
rect 12448 399978 12768 400046
rect 12448 399922 12518 399978
rect 12574 399922 12642 399978
rect 12698 399922 12768 399978
rect 12448 399888 12768 399922
rect 43168 400350 43488 400384
rect 43168 400294 43238 400350
rect 43294 400294 43362 400350
rect 43418 400294 43488 400350
rect 43168 400226 43488 400294
rect 43168 400170 43238 400226
rect 43294 400170 43362 400226
rect 43418 400170 43488 400226
rect 43168 400102 43488 400170
rect 43168 400046 43238 400102
rect 43294 400046 43362 400102
rect 43418 400046 43488 400102
rect 43168 399978 43488 400046
rect 43168 399922 43238 399978
rect 43294 399922 43362 399978
rect 43418 399922 43488 399978
rect 43168 399888 43488 399922
rect 73888 400350 74208 400384
rect 73888 400294 73958 400350
rect 74014 400294 74082 400350
rect 74138 400294 74208 400350
rect 73888 400226 74208 400294
rect 73888 400170 73958 400226
rect 74014 400170 74082 400226
rect 74138 400170 74208 400226
rect 73888 400102 74208 400170
rect 73888 400046 73958 400102
rect 74014 400046 74082 400102
rect 74138 400046 74208 400102
rect 73888 399978 74208 400046
rect 73888 399922 73958 399978
rect 74014 399922 74082 399978
rect 74138 399922 74208 399978
rect 73888 399888 74208 399922
rect 104608 400350 104928 400384
rect 104608 400294 104678 400350
rect 104734 400294 104802 400350
rect 104858 400294 104928 400350
rect 104608 400226 104928 400294
rect 104608 400170 104678 400226
rect 104734 400170 104802 400226
rect 104858 400170 104928 400226
rect 104608 400102 104928 400170
rect 104608 400046 104678 400102
rect 104734 400046 104802 400102
rect 104858 400046 104928 400102
rect 104608 399978 104928 400046
rect 104608 399922 104678 399978
rect 104734 399922 104802 399978
rect 104858 399922 104928 399978
rect 104608 399888 104928 399922
rect 135328 400350 135648 400384
rect 135328 400294 135398 400350
rect 135454 400294 135522 400350
rect 135578 400294 135648 400350
rect 135328 400226 135648 400294
rect 135328 400170 135398 400226
rect 135454 400170 135522 400226
rect 135578 400170 135648 400226
rect 135328 400102 135648 400170
rect 135328 400046 135398 400102
rect 135454 400046 135522 400102
rect 135578 400046 135648 400102
rect 135328 399978 135648 400046
rect 135328 399922 135398 399978
rect 135454 399922 135522 399978
rect 135578 399922 135648 399978
rect 135328 399888 135648 399922
rect 166048 400350 166368 400384
rect 166048 400294 166118 400350
rect 166174 400294 166242 400350
rect 166298 400294 166368 400350
rect 166048 400226 166368 400294
rect 166048 400170 166118 400226
rect 166174 400170 166242 400226
rect 166298 400170 166368 400226
rect 166048 400102 166368 400170
rect 166048 400046 166118 400102
rect 166174 400046 166242 400102
rect 166298 400046 166368 400102
rect 166048 399978 166368 400046
rect 166048 399922 166118 399978
rect 166174 399922 166242 399978
rect 166298 399922 166368 399978
rect 166048 399888 166368 399922
rect 196768 400350 197088 400384
rect 196768 400294 196838 400350
rect 196894 400294 196962 400350
rect 197018 400294 197088 400350
rect 196768 400226 197088 400294
rect 196768 400170 196838 400226
rect 196894 400170 196962 400226
rect 197018 400170 197088 400226
rect 196768 400102 197088 400170
rect 196768 400046 196838 400102
rect 196894 400046 196962 400102
rect 197018 400046 197088 400102
rect 196768 399978 197088 400046
rect 196768 399922 196838 399978
rect 196894 399922 196962 399978
rect 197018 399922 197088 399978
rect 196768 399888 197088 399922
rect 227488 400350 227808 400384
rect 227488 400294 227558 400350
rect 227614 400294 227682 400350
rect 227738 400294 227808 400350
rect 227488 400226 227808 400294
rect 227488 400170 227558 400226
rect 227614 400170 227682 400226
rect 227738 400170 227808 400226
rect 227488 400102 227808 400170
rect 227488 400046 227558 400102
rect 227614 400046 227682 400102
rect 227738 400046 227808 400102
rect 227488 399978 227808 400046
rect 227488 399922 227558 399978
rect 227614 399922 227682 399978
rect 227738 399922 227808 399978
rect 227488 399888 227808 399922
rect 258208 400350 258528 400384
rect 258208 400294 258278 400350
rect 258334 400294 258402 400350
rect 258458 400294 258528 400350
rect 258208 400226 258528 400294
rect 258208 400170 258278 400226
rect 258334 400170 258402 400226
rect 258458 400170 258528 400226
rect 258208 400102 258528 400170
rect 258208 400046 258278 400102
rect 258334 400046 258402 400102
rect 258458 400046 258528 400102
rect 258208 399978 258528 400046
rect 258208 399922 258278 399978
rect 258334 399922 258402 399978
rect 258458 399922 258528 399978
rect 258208 399888 258528 399922
rect 288928 400350 289248 400384
rect 288928 400294 288998 400350
rect 289054 400294 289122 400350
rect 289178 400294 289248 400350
rect 288928 400226 289248 400294
rect 288928 400170 288998 400226
rect 289054 400170 289122 400226
rect 289178 400170 289248 400226
rect 288928 400102 289248 400170
rect 288928 400046 288998 400102
rect 289054 400046 289122 400102
rect 289178 400046 289248 400102
rect 288928 399978 289248 400046
rect 288928 399922 288998 399978
rect 289054 399922 289122 399978
rect 289178 399922 289248 399978
rect 288928 399888 289248 399922
rect 319648 400350 319968 400384
rect 319648 400294 319718 400350
rect 319774 400294 319842 400350
rect 319898 400294 319968 400350
rect 319648 400226 319968 400294
rect 319648 400170 319718 400226
rect 319774 400170 319842 400226
rect 319898 400170 319968 400226
rect 319648 400102 319968 400170
rect 319648 400046 319718 400102
rect 319774 400046 319842 400102
rect 319898 400046 319968 400102
rect 319648 399978 319968 400046
rect 319648 399922 319718 399978
rect 319774 399922 319842 399978
rect 319898 399922 319968 399978
rect 319648 399888 319968 399922
rect 350368 400350 350688 400384
rect 350368 400294 350438 400350
rect 350494 400294 350562 400350
rect 350618 400294 350688 400350
rect 350368 400226 350688 400294
rect 350368 400170 350438 400226
rect 350494 400170 350562 400226
rect 350618 400170 350688 400226
rect 350368 400102 350688 400170
rect 350368 400046 350438 400102
rect 350494 400046 350562 400102
rect 350618 400046 350688 400102
rect 350368 399978 350688 400046
rect 350368 399922 350438 399978
rect 350494 399922 350562 399978
rect 350618 399922 350688 399978
rect 350368 399888 350688 399922
rect 381088 400350 381408 400384
rect 381088 400294 381158 400350
rect 381214 400294 381282 400350
rect 381338 400294 381408 400350
rect 381088 400226 381408 400294
rect 381088 400170 381158 400226
rect 381214 400170 381282 400226
rect 381338 400170 381408 400226
rect 381088 400102 381408 400170
rect 381088 400046 381158 400102
rect 381214 400046 381282 400102
rect 381338 400046 381408 400102
rect 381088 399978 381408 400046
rect 381088 399922 381158 399978
rect 381214 399922 381282 399978
rect 381338 399922 381408 399978
rect 381088 399888 381408 399922
rect 411808 400350 412128 400384
rect 411808 400294 411878 400350
rect 411934 400294 412002 400350
rect 412058 400294 412128 400350
rect 411808 400226 412128 400294
rect 411808 400170 411878 400226
rect 411934 400170 412002 400226
rect 412058 400170 412128 400226
rect 411808 400102 412128 400170
rect 411808 400046 411878 400102
rect 411934 400046 412002 400102
rect 412058 400046 412128 400102
rect 411808 399978 412128 400046
rect 411808 399922 411878 399978
rect 411934 399922 412002 399978
rect 412058 399922 412128 399978
rect 411808 399888 412128 399922
rect 442528 400350 442848 400384
rect 442528 400294 442598 400350
rect 442654 400294 442722 400350
rect 442778 400294 442848 400350
rect 442528 400226 442848 400294
rect 442528 400170 442598 400226
rect 442654 400170 442722 400226
rect 442778 400170 442848 400226
rect 442528 400102 442848 400170
rect 442528 400046 442598 400102
rect 442654 400046 442722 400102
rect 442778 400046 442848 400102
rect 442528 399978 442848 400046
rect 442528 399922 442598 399978
rect 442654 399922 442722 399978
rect 442778 399922 442848 399978
rect 442528 399888 442848 399922
rect 473248 400350 473568 400384
rect 473248 400294 473318 400350
rect 473374 400294 473442 400350
rect 473498 400294 473568 400350
rect 473248 400226 473568 400294
rect 473248 400170 473318 400226
rect 473374 400170 473442 400226
rect 473498 400170 473568 400226
rect 473248 400102 473568 400170
rect 473248 400046 473318 400102
rect 473374 400046 473442 400102
rect 473498 400046 473568 400102
rect 473248 399978 473568 400046
rect 473248 399922 473318 399978
rect 473374 399922 473442 399978
rect 473498 399922 473568 399978
rect 473248 399888 473568 399922
rect 503968 400350 504288 400384
rect 503968 400294 504038 400350
rect 504094 400294 504162 400350
rect 504218 400294 504288 400350
rect 503968 400226 504288 400294
rect 503968 400170 504038 400226
rect 504094 400170 504162 400226
rect 504218 400170 504288 400226
rect 503968 400102 504288 400170
rect 503968 400046 504038 400102
rect 504094 400046 504162 400102
rect 504218 400046 504288 400102
rect 503968 399978 504288 400046
rect 503968 399922 504038 399978
rect 504094 399922 504162 399978
rect 504218 399922 504288 399978
rect 503968 399888 504288 399922
rect 534688 400350 535008 400384
rect 534688 400294 534758 400350
rect 534814 400294 534882 400350
rect 534938 400294 535008 400350
rect 534688 400226 535008 400294
rect 534688 400170 534758 400226
rect 534814 400170 534882 400226
rect 534938 400170 535008 400226
rect 534688 400102 535008 400170
rect 534688 400046 534758 400102
rect 534814 400046 534882 400102
rect 534938 400046 535008 400102
rect 534688 399978 535008 400046
rect 534688 399922 534758 399978
rect 534814 399922 534882 399978
rect 534938 399922 535008 399978
rect 534688 399888 535008 399922
rect 565408 400350 565728 400384
rect 565408 400294 565478 400350
rect 565534 400294 565602 400350
rect 565658 400294 565728 400350
rect 565408 400226 565728 400294
rect 565408 400170 565478 400226
rect 565534 400170 565602 400226
rect 565658 400170 565728 400226
rect 565408 400102 565728 400170
rect 565408 400046 565478 400102
rect 565534 400046 565602 400102
rect 565658 400046 565728 400102
rect 565408 399978 565728 400046
rect 565408 399922 565478 399978
rect 565534 399922 565602 399978
rect 565658 399922 565728 399978
rect 565408 399888 565728 399922
rect 6188 396610 6244 396620
rect 585564 393540 585620 416780
rect 585564 393474 585620 393484
rect 585676 403620 585732 403630
rect 585452 390404 585508 390414
rect 5418 382294 5514 382350
rect 5570 382294 5638 382350
rect 5694 382294 5762 382350
rect 5818 382294 5886 382350
rect 5942 382294 6038 382350
rect 5418 382226 6038 382294
rect 5418 382170 5514 382226
rect 5570 382170 5638 382226
rect 5694 382170 5762 382226
rect 5818 382170 5886 382226
rect 5942 382170 6038 382226
rect 5418 382102 6038 382170
rect 5418 382046 5514 382102
rect 5570 382046 5638 382102
rect 5694 382046 5762 382102
rect 5818 382046 5886 382102
rect 5942 382046 6038 382102
rect 5418 381978 6038 382046
rect 5418 381922 5514 381978
rect 5570 381922 5638 381978
rect 5694 381922 5762 381978
rect 5818 381922 5886 381978
rect 5942 381922 6038 381978
rect 5418 364350 6038 381922
rect 6412 389620 6468 389630
rect 6412 375620 6468 389564
rect 27808 388350 28128 388384
rect 27808 388294 27878 388350
rect 27934 388294 28002 388350
rect 28058 388294 28128 388350
rect 27808 388226 28128 388294
rect 27808 388170 27878 388226
rect 27934 388170 28002 388226
rect 28058 388170 28128 388226
rect 27808 388102 28128 388170
rect 27808 388046 27878 388102
rect 27934 388046 28002 388102
rect 28058 388046 28128 388102
rect 27808 387978 28128 388046
rect 27808 387922 27878 387978
rect 27934 387922 28002 387978
rect 28058 387922 28128 387978
rect 27808 387888 28128 387922
rect 58528 388350 58848 388384
rect 58528 388294 58598 388350
rect 58654 388294 58722 388350
rect 58778 388294 58848 388350
rect 58528 388226 58848 388294
rect 58528 388170 58598 388226
rect 58654 388170 58722 388226
rect 58778 388170 58848 388226
rect 58528 388102 58848 388170
rect 58528 388046 58598 388102
rect 58654 388046 58722 388102
rect 58778 388046 58848 388102
rect 58528 387978 58848 388046
rect 58528 387922 58598 387978
rect 58654 387922 58722 387978
rect 58778 387922 58848 387978
rect 58528 387888 58848 387922
rect 89248 388350 89568 388384
rect 89248 388294 89318 388350
rect 89374 388294 89442 388350
rect 89498 388294 89568 388350
rect 89248 388226 89568 388294
rect 89248 388170 89318 388226
rect 89374 388170 89442 388226
rect 89498 388170 89568 388226
rect 89248 388102 89568 388170
rect 89248 388046 89318 388102
rect 89374 388046 89442 388102
rect 89498 388046 89568 388102
rect 89248 387978 89568 388046
rect 89248 387922 89318 387978
rect 89374 387922 89442 387978
rect 89498 387922 89568 387978
rect 89248 387888 89568 387922
rect 119968 388350 120288 388384
rect 119968 388294 120038 388350
rect 120094 388294 120162 388350
rect 120218 388294 120288 388350
rect 119968 388226 120288 388294
rect 119968 388170 120038 388226
rect 120094 388170 120162 388226
rect 120218 388170 120288 388226
rect 119968 388102 120288 388170
rect 119968 388046 120038 388102
rect 120094 388046 120162 388102
rect 120218 388046 120288 388102
rect 119968 387978 120288 388046
rect 119968 387922 120038 387978
rect 120094 387922 120162 387978
rect 120218 387922 120288 387978
rect 119968 387888 120288 387922
rect 150688 388350 151008 388384
rect 150688 388294 150758 388350
rect 150814 388294 150882 388350
rect 150938 388294 151008 388350
rect 150688 388226 151008 388294
rect 150688 388170 150758 388226
rect 150814 388170 150882 388226
rect 150938 388170 151008 388226
rect 150688 388102 151008 388170
rect 150688 388046 150758 388102
rect 150814 388046 150882 388102
rect 150938 388046 151008 388102
rect 150688 387978 151008 388046
rect 150688 387922 150758 387978
rect 150814 387922 150882 387978
rect 150938 387922 151008 387978
rect 150688 387888 151008 387922
rect 181408 388350 181728 388384
rect 181408 388294 181478 388350
rect 181534 388294 181602 388350
rect 181658 388294 181728 388350
rect 181408 388226 181728 388294
rect 181408 388170 181478 388226
rect 181534 388170 181602 388226
rect 181658 388170 181728 388226
rect 181408 388102 181728 388170
rect 181408 388046 181478 388102
rect 181534 388046 181602 388102
rect 181658 388046 181728 388102
rect 181408 387978 181728 388046
rect 181408 387922 181478 387978
rect 181534 387922 181602 387978
rect 181658 387922 181728 387978
rect 181408 387888 181728 387922
rect 212128 388350 212448 388384
rect 212128 388294 212198 388350
rect 212254 388294 212322 388350
rect 212378 388294 212448 388350
rect 212128 388226 212448 388294
rect 212128 388170 212198 388226
rect 212254 388170 212322 388226
rect 212378 388170 212448 388226
rect 212128 388102 212448 388170
rect 212128 388046 212198 388102
rect 212254 388046 212322 388102
rect 212378 388046 212448 388102
rect 212128 387978 212448 388046
rect 212128 387922 212198 387978
rect 212254 387922 212322 387978
rect 212378 387922 212448 387978
rect 212128 387888 212448 387922
rect 242848 388350 243168 388384
rect 242848 388294 242918 388350
rect 242974 388294 243042 388350
rect 243098 388294 243168 388350
rect 242848 388226 243168 388294
rect 242848 388170 242918 388226
rect 242974 388170 243042 388226
rect 243098 388170 243168 388226
rect 242848 388102 243168 388170
rect 242848 388046 242918 388102
rect 242974 388046 243042 388102
rect 243098 388046 243168 388102
rect 242848 387978 243168 388046
rect 242848 387922 242918 387978
rect 242974 387922 243042 387978
rect 243098 387922 243168 387978
rect 242848 387888 243168 387922
rect 273568 388350 273888 388384
rect 273568 388294 273638 388350
rect 273694 388294 273762 388350
rect 273818 388294 273888 388350
rect 273568 388226 273888 388294
rect 273568 388170 273638 388226
rect 273694 388170 273762 388226
rect 273818 388170 273888 388226
rect 273568 388102 273888 388170
rect 273568 388046 273638 388102
rect 273694 388046 273762 388102
rect 273818 388046 273888 388102
rect 273568 387978 273888 388046
rect 273568 387922 273638 387978
rect 273694 387922 273762 387978
rect 273818 387922 273888 387978
rect 273568 387888 273888 387922
rect 304288 388350 304608 388384
rect 304288 388294 304358 388350
rect 304414 388294 304482 388350
rect 304538 388294 304608 388350
rect 304288 388226 304608 388294
rect 304288 388170 304358 388226
rect 304414 388170 304482 388226
rect 304538 388170 304608 388226
rect 304288 388102 304608 388170
rect 304288 388046 304358 388102
rect 304414 388046 304482 388102
rect 304538 388046 304608 388102
rect 304288 387978 304608 388046
rect 304288 387922 304358 387978
rect 304414 387922 304482 387978
rect 304538 387922 304608 387978
rect 304288 387888 304608 387922
rect 335008 388350 335328 388384
rect 335008 388294 335078 388350
rect 335134 388294 335202 388350
rect 335258 388294 335328 388350
rect 335008 388226 335328 388294
rect 335008 388170 335078 388226
rect 335134 388170 335202 388226
rect 335258 388170 335328 388226
rect 335008 388102 335328 388170
rect 335008 388046 335078 388102
rect 335134 388046 335202 388102
rect 335258 388046 335328 388102
rect 335008 387978 335328 388046
rect 335008 387922 335078 387978
rect 335134 387922 335202 387978
rect 335258 387922 335328 387978
rect 335008 387888 335328 387922
rect 365728 388350 366048 388384
rect 365728 388294 365798 388350
rect 365854 388294 365922 388350
rect 365978 388294 366048 388350
rect 365728 388226 366048 388294
rect 365728 388170 365798 388226
rect 365854 388170 365922 388226
rect 365978 388170 366048 388226
rect 365728 388102 366048 388170
rect 365728 388046 365798 388102
rect 365854 388046 365922 388102
rect 365978 388046 366048 388102
rect 365728 387978 366048 388046
rect 365728 387922 365798 387978
rect 365854 387922 365922 387978
rect 365978 387922 366048 387978
rect 365728 387888 366048 387922
rect 396448 388350 396768 388384
rect 396448 388294 396518 388350
rect 396574 388294 396642 388350
rect 396698 388294 396768 388350
rect 396448 388226 396768 388294
rect 396448 388170 396518 388226
rect 396574 388170 396642 388226
rect 396698 388170 396768 388226
rect 396448 388102 396768 388170
rect 396448 388046 396518 388102
rect 396574 388046 396642 388102
rect 396698 388046 396768 388102
rect 396448 387978 396768 388046
rect 396448 387922 396518 387978
rect 396574 387922 396642 387978
rect 396698 387922 396768 387978
rect 396448 387888 396768 387922
rect 427168 388350 427488 388384
rect 427168 388294 427238 388350
rect 427294 388294 427362 388350
rect 427418 388294 427488 388350
rect 427168 388226 427488 388294
rect 427168 388170 427238 388226
rect 427294 388170 427362 388226
rect 427418 388170 427488 388226
rect 427168 388102 427488 388170
rect 427168 388046 427238 388102
rect 427294 388046 427362 388102
rect 427418 388046 427488 388102
rect 427168 387978 427488 388046
rect 427168 387922 427238 387978
rect 427294 387922 427362 387978
rect 427418 387922 427488 387978
rect 427168 387888 427488 387922
rect 457888 388350 458208 388384
rect 457888 388294 457958 388350
rect 458014 388294 458082 388350
rect 458138 388294 458208 388350
rect 457888 388226 458208 388294
rect 457888 388170 457958 388226
rect 458014 388170 458082 388226
rect 458138 388170 458208 388226
rect 457888 388102 458208 388170
rect 457888 388046 457958 388102
rect 458014 388046 458082 388102
rect 458138 388046 458208 388102
rect 457888 387978 458208 388046
rect 457888 387922 457958 387978
rect 458014 387922 458082 387978
rect 458138 387922 458208 387978
rect 457888 387888 458208 387922
rect 488608 388350 488928 388384
rect 488608 388294 488678 388350
rect 488734 388294 488802 388350
rect 488858 388294 488928 388350
rect 488608 388226 488928 388294
rect 488608 388170 488678 388226
rect 488734 388170 488802 388226
rect 488858 388170 488928 388226
rect 488608 388102 488928 388170
rect 488608 388046 488678 388102
rect 488734 388046 488802 388102
rect 488858 388046 488928 388102
rect 488608 387978 488928 388046
rect 488608 387922 488678 387978
rect 488734 387922 488802 387978
rect 488858 387922 488928 387978
rect 488608 387888 488928 387922
rect 519328 388350 519648 388384
rect 519328 388294 519398 388350
rect 519454 388294 519522 388350
rect 519578 388294 519648 388350
rect 519328 388226 519648 388294
rect 519328 388170 519398 388226
rect 519454 388170 519522 388226
rect 519578 388170 519648 388226
rect 519328 388102 519648 388170
rect 519328 388046 519398 388102
rect 519454 388046 519522 388102
rect 519578 388046 519648 388102
rect 519328 387978 519648 388046
rect 519328 387922 519398 387978
rect 519454 387922 519522 387978
rect 519578 387922 519648 387978
rect 519328 387888 519648 387922
rect 550048 388350 550368 388384
rect 550048 388294 550118 388350
rect 550174 388294 550242 388350
rect 550298 388294 550368 388350
rect 550048 388226 550368 388294
rect 550048 388170 550118 388226
rect 550174 388170 550242 388226
rect 550298 388170 550368 388226
rect 550048 388102 550368 388170
rect 550048 388046 550118 388102
rect 550174 388046 550242 388102
rect 550298 388046 550368 388102
rect 550048 387978 550368 388046
rect 550048 387922 550118 387978
rect 550174 387922 550242 387978
rect 550298 387922 550368 387978
rect 550048 387888 550368 387922
rect 12448 382350 12768 382384
rect 12448 382294 12518 382350
rect 12574 382294 12642 382350
rect 12698 382294 12768 382350
rect 12448 382226 12768 382294
rect 12448 382170 12518 382226
rect 12574 382170 12642 382226
rect 12698 382170 12768 382226
rect 12448 382102 12768 382170
rect 12448 382046 12518 382102
rect 12574 382046 12642 382102
rect 12698 382046 12768 382102
rect 12448 381978 12768 382046
rect 12448 381922 12518 381978
rect 12574 381922 12642 381978
rect 12698 381922 12768 381978
rect 12448 381888 12768 381922
rect 43168 382350 43488 382384
rect 43168 382294 43238 382350
rect 43294 382294 43362 382350
rect 43418 382294 43488 382350
rect 43168 382226 43488 382294
rect 43168 382170 43238 382226
rect 43294 382170 43362 382226
rect 43418 382170 43488 382226
rect 43168 382102 43488 382170
rect 43168 382046 43238 382102
rect 43294 382046 43362 382102
rect 43418 382046 43488 382102
rect 43168 381978 43488 382046
rect 43168 381922 43238 381978
rect 43294 381922 43362 381978
rect 43418 381922 43488 381978
rect 43168 381888 43488 381922
rect 73888 382350 74208 382384
rect 73888 382294 73958 382350
rect 74014 382294 74082 382350
rect 74138 382294 74208 382350
rect 73888 382226 74208 382294
rect 73888 382170 73958 382226
rect 74014 382170 74082 382226
rect 74138 382170 74208 382226
rect 73888 382102 74208 382170
rect 73888 382046 73958 382102
rect 74014 382046 74082 382102
rect 74138 382046 74208 382102
rect 73888 381978 74208 382046
rect 73888 381922 73958 381978
rect 74014 381922 74082 381978
rect 74138 381922 74208 381978
rect 73888 381888 74208 381922
rect 104608 382350 104928 382384
rect 104608 382294 104678 382350
rect 104734 382294 104802 382350
rect 104858 382294 104928 382350
rect 104608 382226 104928 382294
rect 104608 382170 104678 382226
rect 104734 382170 104802 382226
rect 104858 382170 104928 382226
rect 104608 382102 104928 382170
rect 104608 382046 104678 382102
rect 104734 382046 104802 382102
rect 104858 382046 104928 382102
rect 104608 381978 104928 382046
rect 104608 381922 104678 381978
rect 104734 381922 104802 381978
rect 104858 381922 104928 381978
rect 104608 381888 104928 381922
rect 135328 382350 135648 382384
rect 135328 382294 135398 382350
rect 135454 382294 135522 382350
rect 135578 382294 135648 382350
rect 135328 382226 135648 382294
rect 135328 382170 135398 382226
rect 135454 382170 135522 382226
rect 135578 382170 135648 382226
rect 135328 382102 135648 382170
rect 135328 382046 135398 382102
rect 135454 382046 135522 382102
rect 135578 382046 135648 382102
rect 135328 381978 135648 382046
rect 135328 381922 135398 381978
rect 135454 381922 135522 381978
rect 135578 381922 135648 381978
rect 135328 381888 135648 381922
rect 166048 382350 166368 382384
rect 166048 382294 166118 382350
rect 166174 382294 166242 382350
rect 166298 382294 166368 382350
rect 166048 382226 166368 382294
rect 166048 382170 166118 382226
rect 166174 382170 166242 382226
rect 166298 382170 166368 382226
rect 166048 382102 166368 382170
rect 166048 382046 166118 382102
rect 166174 382046 166242 382102
rect 166298 382046 166368 382102
rect 166048 381978 166368 382046
rect 166048 381922 166118 381978
rect 166174 381922 166242 381978
rect 166298 381922 166368 381978
rect 166048 381888 166368 381922
rect 196768 382350 197088 382384
rect 196768 382294 196838 382350
rect 196894 382294 196962 382350
rect 197018 382294 197088 382350
rect 196768 382226 197088 382294
rect 196768 382170 196838 382226
rect 196894 382170 196962 382226
rect 197018 382170 197088 382226
rect 196768 382102 197088 382170
rect 196768 382046 196838 382102
rect 196894 382046 196962 382102
rect 197018 382046 197088 382102
rect 196768 381978 197088 382046
rect 196768 381922 196838 381978
rect 196894 381922 196962 381978
rect 197018 381922 197088 381978
rect 196768 381888 197088 381922
rect 227488 382350 227808 382384
rect 227488 382294 227558 382350
rect 227614 382294 227682 382350
rect 227738 382294 227808 382350
rect 227488 382226 227808 382294
rect 227488 382170 227558 382226
rect 227614 382170 227682 382226
rect 227738 382170 227808 382226
rect 227488 382102 227808 382170
rect 227488 382046 227558 382102
rect 227614 382046 227682 382102
rect 227738 382046 227808 382102
rect 227488 381978 227808 382046
rect 227488 381922 227558 381978
rect 227614 381922 227682 381978
rect 227738 381922 227808 381978
rect 227488 381888 227808 381922
rect 258208 382350 258528 382384
rect 258208 382294 258278 382350
rect 258334 382294 258402 382350
rect 258458 382294 258528 382350
rect 258208 382226 258528 382294
rect 258208 382170 258278 382226
rect 258334 382170 258402 382226
rect 258458 382170 258528 382226
rect 258208 382102 258528 382170
rect 258208 382046 258278 382102
rect 258334 382046 258402 382102
rect 258458 382046 258528 382102
rect 258208 381978 258528 382046
rect 258208 381922 258278 381978
rect 258334 381922 258402 381978
rect 258458 381922 258528 381978
rect 258208 381888 258528 381922
rect 288928 382350 289248 382384
rect 288928 382294 288998 382350
rect 289054 382294 289122 382350
rect 289178 382294 289248 382350
rect 288928 382226 289248 382294
rect 288928 382170 288998 382226
rect 289054 382170 289122 382226
rect 289178 382170 289248 382226
rect 288928 382102 289248 382170
rect 288928 382046 288998 382102
rect 289054 382046 289122 382102
rect 289178 382046 289248 382102
rect 288928 381978 289248 382046
rect 288928 381922 288998 381978
rect 289054 381922 289122 381978
rect 289178 381922 289248 381978
rect 288928 381888 289248 381922
rect 319648 382350 319968 382384
rect 319648 382294 319718 382350
rect 319774 382294 319842 382350
rect 319898 382294 319968 382350
rect 319648 382226 319968 382294
rect 319648 382170 319718 382226
rect 319774 382170 319842 382226
rect 319898 382170 319968 382226
rect 319648 382102 319968 382170
rect 319648 382046 319718 382102
rect 319774 382046 319842 382102
rect 319898 382046 319968 382102
rect 319648 381978 319968 382046
rect 319648 381922 319718 381978
rect 319774 381922 319842 381978
rect 319898 381922 319968 381978
rect 319648 381888 319968 381922
rect 350368 382350 350688 382384
rect 350368 382294 350438 382350
rect 350494 382294 350562 382350
rect 350618 382294 350688 382350
rect 350368 382226 350688 382294
rect 350368 382170 350438 382226
rect 350494 382170 350562 382226
rect 350618 382170 350688 382226
rect 350368 382102 350688 382170
rect 350368 382046 350438 382102
rect 350494 382046 350562 382102
rect 350618 382046 350688 382102
rect 350368 381978 350688 382046
rect 350368 381922 350438 381978
rect 350494 381922 350562 381978
rect 350618 381922 350688 381978
rect 350368 381888 350688 381922
rect 381088 382350 381408 382384
rect 381088 382294 381158 382350
rect 381214 382294 381282 382350
rect 381338 382294 381408 382350
rect 381088 382226 381408 382294
rect 381088 382170 381158 382226
rect 381214 382170 381282 382226
rect 381338 382170 381408 382226
rect 381088 382102 381408 382170
rect 381088 382046 381158 382102
rect 381214 382046 381282 382102
rect 381338 382046 381408 382102
rect 381088 381978 381408 382046
rect 381088 381922 381158 381978
rect 381214 381922 381282 381978
rect 381338 381922 381408 381978
rect 381088 381888 381408 381922
rect 411808 382350 412128 382384
rect 411808 382294 411878 382350
rect 411934 382294 412002 382350
rect 412058 382294 412128 382350
rect 411808 382226 412128 382294
rect 411808 382170 411878 382226
rect 411934 382170 412002 382226
rect 412058 382170 412128 382226
rect 411808 382102 412128 382170
rect 411808 382046 411878 382102
rect 411934 382046 412002 382102
rect 412058 382046 412128 382102
rect 411808 381978 412128 382046
rect 411808 381922 411878 381978
rect 411934 381922 412002 381978
rect 412058 381922 412128 381978
rect 411808 381888 412128 381922
rect 442528 382350 442848 382384
rect 442528 382294 442598 382350
rect 442654 382294 442722 382350
rect 442778 382294 442848 382350
rect 442528 382226 442848 382294
rect 442528 382170 442598 382226
rect 442654 382170 442722 382226
rect 442778 382170 442848 382226
rect 442528 382102 442848 382170
rect 442528 382046 442598 382102
rect 442654 382046 442722 382102
rect 442778 382046 442848 382102
rect 442528 381978 442848 382046
rect 442528 381922 442598 381978
rect 442654 381922 442722 381978
rect 442778 381922 442848 381978
rect 442528 381888 442848 381922
rect 473248 382350 473568 382384
rect 473248 382294 473318 382350
rect 473374 382294 473442 382350
rect 473498 382294 473568 382350
rect 473248 382226 473568 382294
rect 473248 382170 473318 382226
rect 473374 382170 473442 382226
rect 473498 382170 473568 382226
rect 473248 382102 473568 382170
rect 473248 382046 473318 382102
rect 473374 382046 473442 382102
rect 473498 382046 473568 382102
rect 473248 381978 473568 382046
rect 473248 381922 473318 381978
rect 473374 381922 473442 381978
rect 473498 381922 473568 381978
rect 473248 381888 473568 381922
rect 503968 382350 504288 382384
rect 503968 382294 504038 382350
rect 504094 382294 504162 382350
rect 504218 382294 504288 382350
rect 503968 382226 504288 382294
rect 503968 382170 504038 382226
rect 504094 382170 504162 382226
rect 504218 382170 504288 382226
rect 503968 382102 504288 382170
rect 503968 382046 504038 382102
rect 504094 382046 504162 382102
rect 504218 382046 504288 382102
rect 503968 381978 504288 382046
rect 503968 381922 504038 381978
rect 504094 381922 504162 381978
rect 504218 381922 504288 381978
rect 503968 381888 504288 381922
rect 534688 382350 535008 382384
rect 534688 382294 534758 382350
rect 534814 382294 534882 382350
rect 534938 382294 535008 382350
rect 534688 382226 535008 382294
rect 534688 382170 534758 382226
rect 534814 382170 534882 382226
rect 534938 382170 535008 382226
rect 534688 382102 535008 382170
rect 534688 382046 534758 382102
rect 534814 382046 534882 382102
rect 534938 382046 535008 382102
rect 534688 381978 535008 382046
rect 534688 381922 534758 381978
rect 534814 381922 534882 381978
rect 534938 381922 535008 381978
rect 534688 381888 535008 381922
rect 565408 382350 565728 382384
rect 565408 382294 565478 382350
rect 565534 382294 565602 382350
rect 565658 382294 565728 382350
rect 565408 382226 565728 382294
rect 565408 382170 565478 382226
rect 565534 382170 565602 382226
rect 565658 382170 565728 382226
rect 565408 382102 565728 382170
rect 565408 382046 565478 382102
rect 565534 382046 565602 382102
rect 565658 382046 565728 382102
rect 565408 381978 565728 382046
rect 565408 381922 565478 381978
rect 565534 381922 565602 381978
rect 565658 381922 565728 381978
rect 565408 381888 565728 381922
rect 6412 375554 6468 375564
rect 5418 364294 5514 364350
rect 5570 364294 5638 364350
rect 5694 364294 5762 364350
rect 5818 364294 5886 364350
rect 5942 364294 6038 364350
rect 5418 364226 6038 364294
rect 5418 364170 5514 364226
rect 5570 364170 5638 364226
rect 5694 364170 5762 364226
rect 5818 364170 5886 364226
rect 5942 364170 6038 364226
rect 5418 364102 6038 364170
rect 5418 364046 5514 364102
rect 5570 364046 5638 364102
rect 5694 364046 5762 364102
rect 5818 364046 5886 364102
rect 5942 364046 6038 364102
rect 5418 363978 6038 364046
rect 5418 363922 5514 363978
rect 5570 363922 5638 363978
rect 5694 363922 5762 363978
rect 5818 363922 5886 363978
rect 5942 363922 6038 363978
rect -956 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 -336 346350
rect -956 346226 -336 346294
rect -956 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 -336 346226
rect -956 346102 -336 346170
rect -956 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 -336 346102
rect -956 345978 -336 346046
rect -956 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 -336 345978
rect -956 328350 -336 345922
rect 4172 361396 4228 361406
rect 4172 344036 4228 361340
rect 4172 343970 4228 343980
rect 5418 346350 6038 363922
rect 6188 375508 6244 375518
rect 6188 354564 6244 375452
rect 27808 370350 28128 370384
rect 27808 370294 27878 370350
rect 27934 370294 28002 370350
rect 28058 370294 28128 370350
rect 27808 370226 28128 370294
rect 27808 370170 27878 370226
rect 27934 370170 28002 370226
rect 28058 370170 28128 370226
rect 27808 370102 28128 370170
rect 27808 370046 27878 370102
rect 27934 370046 28002 370102
rect 28058 370046 28128 370102
rect 27808 369978 28128 370046
rect 27808 369922 27878 369978
rect 27934 369922 28002 369978
rect 28058 369922 28128 369978
rect 27808 369888 28128 369922
rect 58528 370350 58848 370384
rect 58528 370294 58598 370350
rect 58654 370294 58722 370350
rect 58778 370294 58848 370350
rect 58528 370226 58848 370294
rect 58528 370170 58598 370226
rect 58654 370170 58722 370226
rect 58778 370170 58848 370226
rect 58528 370102 58848 370170
rect 58528 370046 58598 370102
rect 58654 370046 58722 370102
rect 58778 370046 58848 370102
rect 58528 369978 58848 370046
rect 58528 369922 58598 369978
rect 58654 369922 58722 369978
rect 58778 369922 58848 369978
rect 58528 369888 58848 369922
rect 89248 370350 89568 370384
rect 89248 370294 89318 370350
rect 89374 370294 89442 370350
rect 89498 370294 89568 370350
rect 89248 370226 89568 370294
rect 89248 370170 89318 370226
rect 89374 370170 89442 370226
rect 89498 370170 89568 370226
rect 89248 370102 89568 370170
rect 89248 370046 89318 370102
rect 89374 370046 89442 370102
rect 89498 370046 89568 370102
rect 89248 369978 89568 370046
rect 89248 369922 89318 369978
rect 89374 369922 89442 369978
rect 89498 369922 89568 369978
rect 89248 369888 89568 369922
rect 119968 370350 120288 370384
rect 119968 370294 120038 370350
rect 120094 370294 120162 370350
rect 120218 370294 120288 370350
rect 119968 370226 120288 370294
rect 119968 370170 120038 370226
rect 120094 370170 120162 370226
rect 120218 370170 120288 370226
rect 119968 370102 120288 370170
rect 119968 370046 120038 370102
rect 120094 370046 120162 370102
rect 120218 370046 120288 370102
rect 119968 369978 120288 370046
rect 119968 369922 120038 369978
rect 120094 369922 120162 369978
rect 120218 369922 120288 369978
rect 119968 369888 120288 369922
rect 150688 370350 151008 370384
rect 150688 370294 150758 370350
rect 150814 370294 150882 370350
rect 150938 370294 151008 370350
rect 150688 370226 151008 370294
rect 150688 370170 150758 370226
rect 150814 370170 150882 370226
rect 150938 370170 151008 370226
rect 150688 370102 151008 370170
rect 150688 370046 150758 370102
rect 150814 370046 150882 370102
rect 150938 370046 151008 370102
rect 150688 369978 151008 370046
rect 150688 369922 150758 369978
rect 150814 369922 150882 369978
rect 150938 369922 151008 369978
rect 150688 369888 151008 369922
rect 181408 370350 181728 370384
rect 181408 370294 181478 370350
rect 181534 370294 181602 370350
rect 181658 370294 181728 370350
rect 181408 370226 181728 370294
rect 181408 370170 181478 370226
rect 181534 370170 181602 370226
rect 181658 370170 181728 370226
rect 181408 370102 181728 370170
rect 181408 370046 181478 370102
rect 181534 370046 181602 370102
rect 181658 370046 181728 370102
rect 181408 369978 181728 370046
rect 181408 369922 181478 369978
rect 181534 369922 181602 369978
rect 181658 369922 181728 369978
rect 181408 369888 181728 369922
rect 212128 370350 212448 370384
rect 212128 370294 212198 370350
rect 212254 370294 212322 370350
rect 212378 370294 212448 370350
rect 212128 370226 212448 370294
rect 212128 370170 212198 370226
rect 212254 370170 212322 370226
rect 212378 370170 212448 370226
rect 212128 370102 212448 370170
rect 212128 370046 212198 370102
rect 212254 370046 212322 370102
rect 212378 370046 212448 370102
rect 212128 369978 212448 370046
rect 212128 369922 212198 369978
rect 212254 369922 212322 369978
rect 212378 369922 212448 369978
rect 212128 369888 212448 369922
rect 242848 370350 243168 370384
rect 242848 370294 242918 370350
rect 242974 370294 243042 370350
rect 243098 370294 243168 370350
rect 242848 370226 243168 370294
rect 242848 370170 242918 370226
rect 242974 370170 243042 370226
rect 243098 370170 243168 370226
rect 242848 370102 243168 370170
rect 242848 370046 242918 370102
rect 242974 370046 243042 370102
rect 243098 370046 243168 370102
rect 242848 369978 243168 370046
rect 242848 369922 242918 369978
rect 242974 369922 243042 369978
rect 243098 369922 243168 369978
rect 242848 369888 243168 369922
rect 273568 370350 273888 370384
rect 273568 370294 273638 370350
rect 273694 370294 273762 370350
rect 273818 370294 273888 370350
rect 273568 370226 273888 370294
rect 273568 370170 273638 370226
rect 273694 370170 273762 370226
rect 273818 370170 273888 370226
rect 273568 370102 273888 370170
rect 273568 370046 273638 370102
rect 273694 370046 273762 370102
rect 273818 370046 273888 370102
rect 273568 369978 273888 370046
rect 273568 369922 273638 369978
rect 273694 369922 273762 369978
rect 273818 369922 273888 369978
rect 273568 369888 273888 369922
rect 304288 370350 304608 370384
rect 304288 370294 304358 370350
rect 304414 370294 304482 370350
rect 304538 370294 304608 370350
rect 304288 370226 304608 370294
rect 304288 370170 304358 370226
rect 304414 370170 304482 370226
rect 304538 370170 304608 370226
rect 304288 370102 304608 370170
rect 304288 370046 304358 370102
rect 304414 370046 304482 370102
rect 304538 370046 304608 370102
rect 304288 369978 304608 370046
rect 304288 369922 304358 369978
rect 304414 369922 304482 369978
rect 304538 369922 304608 369978
rect 304288 369888 304608 369922
rect 335008 370350 335328 370384
rect 335008 370294 335078 370350
rect 335134 370294 335202 370350
rect 335258 370294 335328 370350
rect 335008 370226 335328 370294
rect 335008 370170 335078 370226
rect 335134 370170 335202 370226
rect 335258 370170 335328 370226
rect 335008 370102 335328 370170
rect 335008 370046 335078 370102
rect 335134 370046 335202 370102
rect 335258 370046 335328 370102
rect 335008 369978 335328 370046
rect 335008 369922 335078 369978
rect 335134 369922 335202 369978
rect 335258 369922 335328 369978
rect 335008 369888 335328 369922
rect 365728 370350 366048 370384
rect 365728 370294 365798 370350
rect 365854 370294 365922 370350
rect 365978 370294 366048 370350
rect 365728 370226 366048 370294
rect 365728 370170 365798 370226
rect 365854 370170 365922 370226
rect 365978 370170 366048 370226
rect 365728 370102 366048 370170
rect 365728 370046 365798 370102
rect 365854 370046 365922 370102
rect 365978 370046 366048 370102
rect 365728 369978 366048 370046
rect 365728 369922 365798 369978
rect 365854 369922 365922 369978
rect 365978 369922 366048 369978
rect 365728 369888 366048 369922
rect 396448 370350 396768 370384
rect 396448 370294 396518 370350
rect 396574 370294 396642 370350
rect 396698 370294 396768 370350
rect 396448 370226 396768 370294
rect 396448 370170 396518 370226
rect 396574 370170 396642 370226
rect 396698 370170 396768 370226
rect 396448 370102 396768 370170
rect 396448 370046 396518 370102
rect 396574 370046 396642 370102
rect 396698 370046 396768 370102
rect 396448 369978 396768 370046
rect 396448 369922 396518 369978
rect 396574 369922 396642 369978
rect 396698 369922 396768 369978
rect 396448 369888 396768 369922
rect 427168 370350 427488 370384
rect 427168 370294 427238 370350
rect 427294 370294 427362 370350
rect 427418 370294 427488 370350
rect 427168 370226 427488 370294
rect 427168 370170 427238 370226
rect 427294 370170 427362 370226
rect 427418 370170 427488 370226
rect 427168 370102 427488 370170
rect 427168 370046 427238 370102
rect 427294 370046 427362 370102
rect 427418 370046 427488 370102
rect 427168 369978 427488 370046
rect 427168 369922 427238 369978
rect 427294 369922 427362 369978
rect 427418 369922 427488 369978
rect 427168 369888 427488 369922
rect 457888 370350 458208 370384
rect 457888 370294 457958 370350
rect 458014 370294 458082 370350
rect 458138 370294 458208 370350
rect 457888 370226 458208 370294
rect 457888 370170 457958 370226
rect 458014 370170 458082 370226
rect 458138 370170 458208 370226
rect 457888 370102 458208 370170
rect 457888 370046 457958 370102
rect 458014 370046 458082 370102
rect 458138 370046 458208 370102
rect 457888 369978 458208 370046
rect 457888 369922 457958 369978
rect 458014 369922 458082 369978
rect 458138 369922 458208 369978
rect 457888 369888 458208 369922
rect 488608 370350 488928 370384
rect 488608 370294 488678 370350
rect 488734 370294 488802 370350
rect 488858 370294 488928 370350
rect 488608 370226 488928 370294
rect 488608 370170 488678 370226
rect 488734 370170 488802 370226
rect 488858 370170 488928 370226
rect 488608 370102 488928 370170
rect 488608 370046 488678 370102
rect 488734 370046 488802 370102
rect 488858 370046 488928 370102
rect 488608 369978 488928 370046
rect 488608 369922 488678 369978
rect 488734 369922 488802 369978
rect 488858 369922 488928 369978
rect 488608 369888 488928 369922
rect 519328 370350 519648 370384
rect 519328 370294 519398 370350
rect 519454 370294 519522 370350
rect 519578 370294 519648 370350
rect 519328 370226 519648 370294
rect 519328 370170 519398 370226
rect 519454 370170 519522 370226
rect 519578 370170 519648 370226
rect 519328 370102 519648 370170
rect 519328 370046 519398 370102
rect 519454 370046 519522 370102
rect 519578 370046 519648 370102
rect 519328 369978 519648 370046
rect 519328 369922 519398 369978
rect 519454 369922 519522 369978
rect 519578 369922 519648 369978
rect 519328 369888 519648 369922
rect 550048 370350 550368 370384
rect 550048 370294 550118 370350
rect 550174 370294 550242 370350
rect 550298 370294 550368 370350
rect 550048 370226 550368 370294
rect 550048 370170 550118 370226
rect 550174 370170 550242 370226
rect 550298 370170 550368 370226
rect 550048 370102 550368 370170
rect 550048 370046 550118 370102
rect 550174 370046 550242 370102
rect 550298 370046 550368 370102
rect 550048 369978 550368 370046
rect 550048 369922 550118 369978
rect 550174 369922 550242 369978
rect 550298 369922 550368 369978
rect 550048 369888 550368 369922
rect 12448 364350 12768 364384
rect 12448 364294 12518 364350
rect 12574 364294 12642 364350
rect 12698 364294 12768 364350
rect 12448 364226 12768 364294
rect 12448 364170 12518 364226
rect 12574 364170 12642 364226
rect 12698 364170 12768 364226
rect 12448 364102 12768 364170
rect 12448 364046 12518 364102
rect 12574 364046 12642 364102
rect 12698 364046 12768 364102
rect 12448 363978 12768 364046
rect 12448 363922 12518 363978
rect 12574 363922 12642 363978
rect 12698 363922 12768 363978
rect 12448 363888 12768 363922
rect 43168 364350 43488 364384
rect 43168 364294 43238 364350
rect 43294 364294 43362 364350
rect 43418 364294 43488 364350
rect 43168 364226 43488 364294
rect 43168 364170 43238 364226
rect 43294 364170 43362 364226
rect 43418 364170 43488 364226
rect 43168 364102 43488 364170
rect 43168 364046 43238 364102
rect 43294 364046 43362 364102
rect 43418 364046 43488 364102
rect 43168 363978 43488 364046
rect 43168 363922 43238 363978
rect 43294 363922 43362 363978
rect 43418 363922 43488 363978
rect 43168 363888 43488 363922
rect 73888 364350 74208 364384
rect 73888 364294 73958 364350
rect 74014 364294 74082 364350
rect 74138 364294 74208 364350
rect 73888 364226 74208 364294
rect 73888 364170 73958 364226
rect 74014 364170 74082 364226
rect 74138 364170 74208 364226
rect 73888 364102 74208 364170
rect 73888 364046 73958 364102
rect 74014 364046 74082 364102
rect 74138 364046 74208 364102
rect 73888 363978 74208 364046
rect 73888 363922 73958 363978
rect 74014 363922 74082 363978
rect 74138 363922 74208 363978
rect 73888 363888 74208 363922
rect 104608 364350 104928 364384
rect 104608 364294 104678 364350
rect 104734 364294 104802 364350
rect 104858 364294 104928 364350
rect 104608 364226 104928 364294
rect 104608 364170 104678 364226
rect 104734 364170 104802 364226
rect 104858 364170 104928 364226
rect 104608 364102 104928 364170
rect 104608 364046 104678 364102
rect 104734 364046 104802 364102
rect 104858 364046 104928 364102
rect 104608 363978 104928 364046
rect 104608 363922 104678 363978
rect 104734 363922 104802 363978
rect 104858 363922 104928 363978
rect 104608 363888 104928 363922
rect 135328 364350 135648 364384
rect 135328 364294 135398 364350
rect 135454 364294 135522 364350
rect 135578 364294 135648 364350
rect 135328 364226 135648 364294
rect 135328 364170 135398 364226
rect 135454 364170 135522 364226
rect 135578 364170 135648 364226
rect 135328 364102 135648 364170
rect 135328 364046 135398 364102
rect 135454 364046 135522 364102
rect 135578 364046 135648 364102
rect 135328 363978 135648 364046
rect 135328 363922 135398 363978
rect 135454 363922 135522 363978
rect 135578 363922 135648 363978
rect 135328 363888 135648 363922
rect 166048 364350 166368 364384
rect 166048 364294 166118 364350
rect 166174 364294 166242 364350
rect 166298 364294 166368 364350
rect 166048 364226 166368 364294
rect 166048 364170 166118 364226
rect 166174 364170 166242 364226
rect 166298 364170 166368 364226
rect 166048 364102 166368 364170
rect 166048 364046 166118 364102
rect 166174 364046 166242 364102
rect 166298 364046 166368 364102
rect 166048 363978 166368 364046
rect 166048 363922 166118 363978
rect 166174 363922 166242 363978
rect 166298 363922 166368 363978
rect 166048 363888 166368 363922
rect 196768 364350 197088 364384
rect 196768 364294 196838 364350
rect 196894 364294 196962 364350
rect 197018 364294 197088 364350
rect 196768 364226 197088 364294
rect 196768 364170 196838 364226
rect 196894 364170 196962 364226
rect 197018 364170 197088 364226
rect 196768 364102 197088 364170
rect 196768 364046 196838 364102
rect 196894 364046 196962 364102
rect 197018 364046 197088 364102
rect 196768 363978 197088 364046
rect 196768 363922 196838 363978
rect 196894 363922 196962 363978
rect 197018 363922 197088 363978
rect 196768 363888 197088 363922
rect 227488 364350 227808 364384
rect 227488 364294 227558 364350
rect 227614 364294 227682 364350
rect 227738 364294 227808 364350
rect 227488 364226 227808 364294
rect 227488 364170 227558 364226
rect 227614 364170 227682 364226
rect 227738 364170 227808 364226
rect 227488 364102 227808 364170
rect 227488 364046 227558 364102
rect 227614 364046 227682 364102
rect 227738 364046 227808 364102
rect 227488 363978 227808 364046
rect 227488 363922 227558 363978
rect 227614 363922 227682 363978
rect 227738 363922 227808 363978
rect 227488 363888 227808 363922
rect 258208 364350 258528 364384
rect 258208 364294 258278 364350
rect 258334 364294 258402 364350
rect 258458 364294 258528 364350
rect 258208 364226 258528 364294
rect 258208 364170 258278 364226
rect 258334 364170 258402 364226
rect 258458 364170 258528 364226
rect 258208 364102 258528 364170
rect 258208 364046 258278 364102
rect 258334 364046 258402 364102
rect 258458 364046 258528 364102
rect 258208 363978 258528 364046
rect 258208 363922 258278 363978
rect 258334 363922 258402 363978
rect 258458 363922 258528 363978
rect 258208 363888 258528 363922
rect 288928 364350 289248 364384
rect 288928 364294 288998 364350
rect 289054 364294 289122 364350
rect 289178 364294 289248 364350
rect 288928 364226 289248 364294
rect 288928 364170 288998 364226
rect 289054 364170 289122 364226
rect 289178 364170 289248 364226
rect 288928 364102 289248 364170
rect 288928 364046 288998 364102
rect 289054 364046 289122 364102
rect 289178 364046 289248 364102
rect 288928 363978 289248 364046
rect 288928 363922 288998 363978
rect 289054 363922 289122 363978
rect 289178 363922 289248 363978
rect 288928 363888 289248 363922
rect 319648 364350 319968 364384
rect 319648 364294 319718 364350
rect 319774 364294 319842 364350
rect 319898 364294 319968 364350
rect 319648 364226 319968 364294
rect 319648 364170 319718 364226
rect 319774 364170 319842 364226
rect 319898 364170 319968 364226
rect 319648 364102 319968 364170
rect 319648 364046 319718 364102
rect 319774 364046 319842 364102
rect 319898 364046 319968 364102
rect 319648 363978 319968 364046
rect 319648 363922 319718 363978
rect 319774 363922 319842 363978
rect 319898 363922 319968 363978
rect 319648 363888 319968 363922
rect 350368 364350 350688 364384
rect 350368 364294 350438 364350
rect 350494 364294 350562 364350
rect 350618 364294 350688 364350
rect 350368 364226 350688 364294
rect 350368 364170 350438 364226
rect 350494 364170 350562 364226
rect 350618 364170 350688 364226
rect 350368 364102 350688 364170
rect 350368 364046 350438 364102
rect 350494 364046 350562 364102
rect 350618 364046 350688 364102
rect 350368 363978 350688 364046
rect 350368 363922 350438 363978
rect 350494 363922 350562 363978
rect 350618 363922 350688 363978
rect 350368 363888 350688 363922
rect 381088 364350 381408 364384
rect 381088 364294 381158 364350
rect 381214 364294 381282 364350
rect 381338 364294 381408 364350
rect 381088 364226 381408 364294
rect 381088 364170 381158 364226
rect 381214 364170 381282 364226
rect 381338 364170 381408 364226
rect 381088 364102 381408 364170
rect 381088 364046 381158 364102
rect 381214 364046 381282 364102
rect 381338 364046 381408 364102
rect 381088 363978 381408 364046
rect 381088 363922 381158 363978
rect 381214 363922 381282 363978
rect 381338 363922 381408 363978
rect 381088 363888 381408 363922
rect 411808 364350 412128 364384
rect 411808 364294 411878 364350
rect 411934 364294 412002 364350
rect 412058 364294 412128 364350
rect 411808 364226 412128 364294
rect 411808 364170 411878 364226
rect 411934 364170 412002 364226
rect 412058 364170 412128 364226
rect 411808 364102 412128 364170
rect 411808 364046 411878 364102
rect 411934 364046 412002 364102
rect 412058 364046 412128 364102
rect 411808 363978 412128 364046
rect 411808 363922 411878 363978
rect 411934 363922 412002 363978
rect 412058 363922 412128 363978
rect 411808 363888 412128 363922
rect 442528 364350 442848 364384
rect 442528 364294 442598 364350
rect 442654 364294 442722 364350
rect 442778 364294 442848 364350
rect 442528 364226 442848 364294
rect 442528 364170 442598 364226
rect 442654 364170 442722 364226
rect 442778 364170 442848 364226
rect 442528 364102 442848 364170
rect 442528 364046 442598 364102
rect 442654 364046 442722 364102
rect 442778 364046 442848 364102
rect 442528 363978 442848 364046
rect 442528 363922 442598 363978
rect 442654 363922 442722 363978
rect 442778 363922 442848 363978
rect 442528 363888 442848 363922
rect 473248 364350 473568 364384
rect 473248 364294 473318 364350
rect 473374 364294 473442 364350
rect 473498 364294 473568 364350
rect 473248 364226 473568 364294
rect 473248 364170 473318 364226
rect 473374 364170 473442 364226
rect 473498 364170 473568 364226
rect 473248 364102 473568 364170
rect 473248 364046 473318 364102
rect 473374 364046 473442 364102
rect 473498 364046 473568 364102
rect 473248 363978 473568 364046
rect 473248 363922 473318 363978
rect 473374 363922 473442 363978
rect 473498 363922 473568 363978
rect 473248 363888 473568 363922
rect 503968 364350 504288 364384
rect 503968 364294 504038 364350
rect 504094 364294 504162 364350
rect 504218 364294 504288 364350
rect 503968 364226 504288 364294
rect 503968 364170 504038 364226
rect 504094 364170 504162 364226
rect 504218 364170 504288 364226
rect 503968 364102 504288 364170
rect 503968 364046 504038 364102
rect 504094 364046 504162 364102
rect 504218 364046 504288 364102
rect 503968 363978 504288 364046
rect 503968 363922 504038 363978
rect 504094 363922 504162 363978
rect 504218 363922 504288 363978
rect 503968 363888 504288 363922
rect 534688 364350 535008 364384
rect 534688 364294 534758 364350
rect 534814 364294 534882 364350
rect 534938 364294 535008 364350
rect 534688 364226 535008 364294
rect 534688 364170 534758 364226
rect 534814 364170 534882 364226
rect 534938 364170 535008 364226
rect 534688 364102 535008 364170
rect 534688 364046 534758 364102
rect 534814 364046 534882 364102
rect 534938 364046 535008 364102
rect 534688 363978 535008 364046
rect 534688 363922 534758 363978
rect 534814 363922 534882 363978
rect 534938 363922 535008 363978
rect 534688 363888 535008 363922
rect 565408 364350 565728 364384
rect 565408 364294 565478 364350
rect 565534 364294 565602 364350
rect 565658 364294 565728 364350
rect 565408 364226 565728 364294
rect 565408 364170 565478 364226
rect 565534 364170 565602 364226
rect 565658 364170 565728 364226
rect 565408 364102 565728 364170
rect 565408 364046 565478 364102
rect 565534 364046 565602 364102
rect 565658 364046 565728 364102
rect 565408 363978 565728 364046
rect 565408 363922 565478 363978
rect 565534 363922 565602 363978
rect 565658 363922 565728 363978
rect 565408 363888 565728 363922
rect 585452 361284 585508 390348
rect 585676 382788 585732 403564
rect 585676 382722 585732 382732
rect 589098 400350 589718 417922
rect 589098 400294 589194 400350
rect 589250 400294 589318 400350
rect 589374 400294 589442 400350
rect 589498 400294 589566 400350
rect 589622 400294 589718 400350
rect 589098 400226 589718 400294
rect 589098 400170 589194 400226
rect 589250 400170 589318 400226
rect 589374 400170 589442 400226
rect 589498 400170 589566 400226
rect 589622 400170 589718 400226
rect 589098 400102 589718 400170
rect 589098 400046 589194 400102
rect 589250 400046 589318 400102
rect 589374 400046 589442 400102
rect 589498 400046 589566 400102
rect 589622 400046 589718 400102
rect 589098 399978 589718 400046
rect 589098 399922 589194 399978
rect 589250 399922 589318 399978
rect 589374 399922 589442 399978
rect 589498 399922 589566 399978
rect 589622 399922 589718 399978
rect 589098 382350 589718 399922
rect 589098 382294 589194 382350
rect 589250 382294 589318 382350
rect 589374 382294 589442 382350
rect 589498 382294 589566 382350
rect 589622 382294 589718 382350
rect 589098 382226 589718 382294
rect 589098 382170 589194 382226
rect 589250 382170 589318 382226
rect 589374 382170 589442 382226
rect 589498 382170 589566 382226
rect 589622 382170 589718 382226
rect 589098 382102 589718 382170
rect 589098 382046 589194 382102
rect 589250 382046 589318 382102
rect 589374 382046 589442 382102
rect 589498 382046 589566 382102
rect 589622 382046 589718 382102
rect 589098 381978 589718 382046
rect 589098 381922 589194 381978
rect 589250 381922 589318 381978
rect 589374 381922 589442 381978
rect 589498 381922 589566 381978
rect 589622 381922 589718 381978
rect 585452 361218 585508 361228
rect 585676 377188 585732 377198
rect 6188 354498 6244 354508
rect 27808 352350 28128 352384
rect 27808 352294 27878 352350
rect 27934 352294 28002 352350
rect 28058 352294 28128 352350
rect 27808 352226 28128 352294
rect 27808 352170 27878 352226
rect 27934 352170 28002 352226
rect 28058 352170 28128 352226
rect 27808 352102 28128 352170
rect 27808 352046 27878 352102
rect 27934 352046 28002 352102
rect 28058 352046 28128 352102
rect 27808 351978 28128 352046
rect 27808 351922 27878 351978
rect 27934 351922 28002 351978
rect 28058 351922 28128 351978
rect 27808 351888 28128 351922
rect 58528 352350 58848 352384
rect 58528 352294 58598 352350
rect 58654 352294 58722 352350
rect 58778 352294 58848 352350
rect 58528 352226 58848 352294
rect 58528 352170 58598 352226
rect 58654 352170 58722 352226
rect 58778 352170 58848 352226
rect 58528 352102 58848 352170
rect 58528 352046 58598 352102
rect 58654 352046 58722 352102
rect 58778 352046 58848 352102
rect 58528 351978 58848 352046
rect 58528 351922 58598 351978
rect 58654 351922 58722 351978
rect 58778 351922 58848 351978
rect 58528 351888 58848 351922
rect 89248 352350 89568 352384
rect 89248 352294 89318 352350
rect 89374 352294 89442 352350
rect 89498 352294 89568 352350
rect 89248 352226 89568 352294
rect 89248 352170 89318 352226
rect 89374 352170 89442 352226
rect 89498 352170 89568 352226
rect 89248 352102 89568 352170
rect 89248 352046 89318 352102
rect 89374 352046 89442 352102
rect 89498 352046 89568 352102
rect 89248 351978 89568 352046
rect 89248 351922 89318 351978
rect 89374 351922 89442 351978
rect 89498 351922 89568 351978
rect 89248 351888 89568 351922
rect 119968 352350 120288 352384
rect 119968 352294 120038 352350
rect 120094 352294 120162 352350
rect 120218 352294 120288 352350
rect 119968 352226 120288 352294
rect 119968 352170 120038 352226
rect 120094 352170 120162 352226
rect 120218 352170 120288 352226
rect 119968 352102 120288 352170
rect 119968 352046 120038 352102
rect 120094 352046 120162 352102
rect 120218 352046 120288 352102
rect 119968 351978 120288 352046
rect 119968 351922 120038 351978
rect 120094 351922 120162 351978
rect 120218 351922 120288 351978
rect 119968 351888 120288 351922
rect 150688 352350 151008 352384
rect 150688 352294 150758 352350
rect 150814 352294 150882 352350
rect 150938 352294 151008 352350
rect 150688 352226 151008 352294
rect 150688 352170 150758 352226
rect 150814 352170 150882 352226
rect 150938 352170 151008 352226
rect 150688 352102 151008 352170
rect 150688 352046 150758 352102
rect 150814 352046 150882 352102
rect 150938 352046 151008 352102
rect 150688 351978 151008 352046
rect 150688 351922 150758 351978
rect 150814 351922 150882 351978
rect 150938 351922 151008 351978
rect 150688 351888 151008 351922
rect 181408 352350 181728 352384
rect 181408 352294 181478 352350
rect 181534 352294 181602 352350
rect 181658 352294 181728 352350
rect 181408 352226 181728 352294
rect 181408 352170 181478 352226
rect 181534 352170 181602 352226
rect 181658 352170 181728 352226
rect 181408 352102 181728 352170
rect 181408 352046 181478 352102
rect 181534 352046 181602 352102
rect 181658 352046 181728 352102
rect 181408 351978 181728 352046
rect 181408 351922 181478 351978
rect 181534 351922 181602 351978
rect 181658 351922 181728 351978
rect 181408 351888 181728 351922
rect 212128 352350 212448 352384
rect 212128 352294 212198 352350
rect 212254 352294 212322 352350
rect 212378 352294 212448 352350
rect 212128 352226 212448 352294
rect 212128 352170 212198 352226
rect 212254 352170 212322 352226
rect 212378 352170 212448 352226
rect 212128 352102 212448 352170
rect 212128 352046 212198 352102
rect 212254 352046 212322 352102
rect 212378 352046 212448 352102
rect 212128 351978 212448 352046
rect 212128 351922 212198 351978
rect 212254 351922 212322 351978
rect 212378 351922 212448 351978
rect 212128 351888 212448 351922
rect 242848 352350 243168 352384
rect 242848 352294 242918 352350
rect 242974 352294 243042 352350
rect 243098 352294 243168 352350
rect 242848 352226 243168 352294
rect 242848 352170 242918 352226
rect 242974 352170 243042 352226
rect 243098 352170 243168 352226
rect 242848 352102 243168 352170
rect 242848 352046 242918 352102
rect 242974 352046 243042 352102
rect 243098 352046 243168 352102
rect 242848 351978 243168 352046
rect 242848 351922 242918 351978
rect 242974 351922 243042 351978
rect 243098 351922 243168 351978
rect 242848 351888 243168 351922
rect 273568 352350 273888 352384
rect 273568 352294 273638 352350
rect 273694 352294 273762 352350
rect 273818 352294 273888 352350
rect 273568 352226 273888 352294
rect 273568 352170 273638 352226
rect 273694 352170 273762 352226
rect 273818 352170 273888 352226
rect 273568 352102 273888 352170
rect 273568 352046 273638 352102
rect 273694 352046 273762 352102
rect 273818 352046 273888 352102
rect 273568 351978 273888 352046
rect 273568 351922 273638 351978
rect 273694 351922 273762 351978
rect 273818 351922 273888 351978
rect 273568 351888 273888 351922
rect 304288 352350 304608 352384
rect 304288 352294 304358 352350
rect 304414 352294 304482 352350
rect 304538 352294 304608 352350
rect 304288 352226 304608 352294
rect 304288 352170 304358 352226
rect 304414 352170 304482 352226
rect 304538 352170 304608 352226
rect 304288 352102 304608 352170
rect 304288 352046 304358 352102
rect 304414 352046 304482 352102
rect 304538 352046 304608 352102
rect 304288 351978 304608 352046
rect 304288 351922 304358 351978
rect 304414 351922 304482 351978
rect 304538 351922 304608 351978
rect 304288 351888 304608 351922
rect 335008 352350 335328 352384
rect 335008 352294 335078 352350
rect 335134 352294 335202 352350
rect 335258 352294 335328 352350
rect 335008 352226 335328 352294
rect 335008 352170 335078 352226
rect 335134 352170 335202 352226
rect 335258 352170 335328 352226
rect 335008 352102 335328 352170
rect 335008 352046 335078 352102
rect 335134 352046 335202 352102
rect 335258 352046 335328 352102
rect 335008 351978 335328 352046
rect 335008 351922 335078 351978
rect 335134 351922 335202 351978
rect 335258 351922 335328 351978
rect 335008 351888 335328 351922
rect 365728 352350 366048 352384
rect 365728 352294 365798 352350
rect 365854 352294 365922 352350
rect 365978 352294 366048 352350
rect 365728 352226 366048 352294
rect 365728 352170 365798 352226
rect 365854 352170 365922 352226
rect 365978 352170 366048 352226
rect 365728 352102 366048 352170
rect 365728 352046 365798 352102
rect 365854 352046 365922 352102
rect 365978 352046 366048 352102
rect 365728 351978 366048 352046
rect 365728 351922 365798 351978
rect 365854 351922 365922 351978
rect 365978 351922 366048 351978
rect 365728 351888 366048 351922
rect 396448 352350 396768 352384
rect 396448 352294 396518 352350
rect 396574 352294 396642 352350
rect 396698 352294 396768 352350
rect 396448 352226 396768 352294
rect 396448 352170 396518 352226
rect 396574 352170 396642 352226
rect 396698 352170 396768 352226
rect 396448 352102 396768 352170
rect 396448 352046 396518 352102
rect 396574 352046 396642 352102
rect 396698 352046 396768 352102
rect 396448 351978 396768 352046
rect 396448 351922 396518 351978
rect 396574 351922 396642 351978
rect 396698 351922 396768 351978
rect 396448 351888 396768 351922
rect 427168 352350 427488 352384
rect 427168 352294 427238 352350
rect 427294 352294 427362 352350
rect 427418 352294 427488 352350
rect 427168 352226 427488 352294
rect 427168 352170 427238 352226
rect 427294 352170 427362 352226
rect 427418 352170 427488 352226
rect 427168 352102 427488 352170
rect 427168 352046 427238 352102
rect 427294 352046 427362 352102
rect 427418 352046 427488 352102
rect 427168 351978 427488 352046
rect 427168 351922 427238 351978
rect 427294 351922 427362 351978
rect 427418 351922 427488 351978
rect 427168 351888 427488 351922
rect 457888 352350 458208 352384
rect 457888 352294 457958 352350
rect 458014 352294 458082 352350
rect 458138 352294 458208 352350
rect 457888 352226 458208 352294
rect 457888 352170 457958 352226
rect 458014 352170 458082 352226
rect 458138 352170 458208 352226
rect 457888 352102 458208 352170
rect 457888 352046 457958 352102
rect 458014 352046 458082 352102
rect 458138 352046 458208 352102
rect 457888 351978 458208 352046
rect 457888 351922 457958 351978
rect 458014 351922 458082 351978
rect 458138 351922 458208 351978
rect 457888 351888 458208 351922
rect 488608 352350 488928 352384
rect 488608 352294 488678 352350
rect 488734 352294 488802 352350
rect 488858 352294 488928 352350
rect 488608 352226 488928 352294
rect 488608 352170 488678 352226
rect 488734 352170 488802 352226
rect 488858 352170 488928 352226
rect 488608 352102 488928 352170
rect 488608 352046 488678 352102
rect 488734 352046 488802 352102
rect 488858 352046 488928 352102
rect 488608 351978 488928 352046
rect 488608 351922 488678 351978
rect 488734 351922 488802 351978
rect 488858 351922 488928 351978
rect 488608 351888 488928 351922
rect 519328 352350 519648 352384
rect 519328 352294 519398 352350
rect 519454 352294 519522 352350
rect 519578 352294 519648 352350
rect 519328 352226 519648 352294
rect 519328 352170 519398 352226
rect 519454 352170 519522 352226
rect 519578 352170 519648 352226
rect 519328 352102 519648 352170
rect 519328 352046 519398 352102
rect 519454 352046 519522 352102
rect 519578 352046 519648 352102
rect 519328 351978 519648 352046
rect 519328 351922 519398 351978
rect 519454 351922 519522 351978
rect 519578 351922 519648 351978
rect 519328 351888 519648 351922
rect 550048 352350 550368 352384
rect 550048 352294 550118 352350
rect 550174 352294 550242 352350
rect 550298 352294 550368 352350
rect 550048 352226 550368 352294
rect 550048 352170 550118 352226
rect 550174 352170 550242 352226
rect 550298 352170 550368 352226
rect 550048 352102 550368 352170
rect 550048 352046 550118 352102
rect 550174 352046 550242 352102
rect 550298 352046 550368 352102
rect 550048 351978 550368 352046
rect 550048 351922 550118 351978
rect 550174 351922 550242 351978
rect 550298 351922 550368 351978
rect 550048 351888 550368 351922
rect 585452 350756 585508 350766
rect 5418 346294 5514 346350
rect 5570 346294 5638 346350
rect 5694 346294 5762 346350
rect 5818 346294 5886 346350
rect 5942 346294 6038 346350
rect 5418 346226 6038 346294
rect 5418 346170 5514 346226
rect 5570 346170 5638 346226
rect 5694 346170 5762 346226
rect 5818 346170 5886 346226
rect 5942 346170 6038 346226
rect 5418 346102 6038 346170
rect 5418 346046 5514 346102
rect 5570 346046 5638 346102
rect 5694 346046 5762 346102
rect 5818 346046 5886 346102
rect 5942 346046 6038 346102
rect 5418 345978 6038 346046
rect 5418 345922 5514 345978
rect 5570 345922 5638 345978
rect 5694 345922 5762 345978
rect 5818 345922 5886 345978
rect 5942 345922 6038 345978
rect -956 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 -336 328350
rect -956 328226 -336 328294
rect -956 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 -336 328226
rect -956 328102 -336 328170
rect -956 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 -336 328102
rect -956 327978 -336 328046
rect -956 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 -336 327978
rect -956 310350 -336 327922
rect 4172 333172 4228 333182
rect 4172 312452 4228 333116
rect 5418 328350 6038 345922
rect 6188 347284 6244 347294
rect 6188 333508 6244 347228
rect 12448 346350 12768 346384
rect 12448 346294 12518 346350
rect 12574 346294 12642 346350
rect 12698 346294 12768 346350
rect 12448 346226 12768 346294
rect 12448 346170 12518 346226
rect 12574 346170 12642 346226
rect 12698 346170 12768 346226
rect 12448 346102 12768 346170
rect 12448 346046 12518 346102
rect 12574 346046 12642 346102
rect 12698 346046 12768 346102
rect 12448 345978 12768 346046
rect 12448 345922 12518 345978
rect 12574 345922 12642 345978
rect 12698 345922 12768 345978
rect 12448 345888 12768 345922
rect 43168 346350 43488 346384
rect 43168 346294 43238 346350
rect 43294 346294 43362 346350
rect 43418 346294 43488 346350
rect 43168 346226 43488 346294
rect 43168 346170 43238 346226
rect 43294 346170 43362 346226
rect 43418 346170 43488 346226
rect 43168 346102 43488 346170
rect 43168 346046 43238 346102
rect 43294 346046 43362 346102
rect 43418 346046 43488 346102
rect 43168 345978 43488 346046
rect 43168 345922 43238 345978
rect 43294 345922 43362 345978
rect 43418 345922 43488 345978
rect 43168 345888 43488 345922
rect 73888 346350 74208 346384
rect 73888 346294 73958 346350
rect 74014 346294 74082 346350
rect 74138 346294 74208 346350
rect 73888 346226 74208 346294
rect 73888 346170 73958 346226
rect 74014 346170 74082 346226
rect 74138 346170 74208 346226
rect 73888 346102 74208 346170
rect 73888 346046 73958 346102
rect 74014 346046 74082 346102
rect 74138 346046 74208 346102
rect 73888 345978 74208 346046
rect 73888 345922 73958 345978
rect 74014 345922 74082 345978
rect 74138 345922 74208 345978
rect 73888 345888 74208 345922
rect 104608 346350 104928 346384
rect 104608 346294 104678 346350
rect 104734 346294 104802 346350
rect 104858 346294 104928 346350
rect 104608 346226 104928 346294
rect 104608 346170 104678 346226
rect 104734 346170 104802 346226
rect 104858 346170 104928 346226
rect 104608 346102 104928 346170
rect 104608 346046 104678 346102
rect 104734 346046 104802 346102
rect 104858 346046 104928 346102
rect 104608 345978 104928 346046
rect 104608 345922 104678 345978
rect 104734 345922 104802 345978
rect 104858 345922 104928 345978
rect 104608 345888 104928 345922
rect 135328 346350 135648 346384
rect 135328 346294 135398 346350
rect 135454 346294 135522 346350
rect 135578 346294 135648 346350
rect 135328 346226 135648 346294
rect 135328 346170 135398 346226
rect 135454 346170 135522 346226
rect 135578 346170 135648 346226
rect 135328 346102 135648 346170
rect 135328 346046 135398 346102
rect 135454 346046 135522 346102
rect 135578 346046 135648 346102
rect 135328 345978 135648 346046
rect 135328 345922 135398 345978
rect 135454 345922 135522 345978
rect 135578 345922 135648 345978
rect 135328 345888 135648 345922
rect 166048 346350 166368 346384
rect 166048 346294 166118 346350
rect 166174 346294 166242 346350
rect 166298 346294 166368 346350
rect 166048 346226 166368 346294
rect 166048 346170 166118 346226
rect 166174 346170 166242 346226
rect 166298 346170 166368 346226
rect 166048 346102 166368 346170
rect 166048 346046 166118 346102
rect 166174 346046 166242 346102
rect 166298 346046 166368 346102
rect 166048 345978 166368 346046
rect 166048 345922 166118 345978
rect 166174 345922 166242 345978
rect 166298 345922 166368 345978
rect 166048 345888 166368 345922
rect 196768 346350 197088 346384
rect 196768 346294 196838 346350
rect 196894 346294 196962 346350
rect 197018 346294 197088 346350
rect 196768 346226 197088 346294
rect 196768 346170 196838 346226
rect 196894 346170 196962 346226
rect 197018 346170 197088 346226
rect 196768 346102 197088 346170
rect 196768 346046 196838 346102
rect 196894 346046 196962 346102
rect 197018 346046 197088 346102
rect 196768 345978 197088 346046
rect 196768 345922 196838 345978
rect 196894 345922 196962 345978
rect 197018 345922 197088 345978
rect 196768 345888 197088 345922
rect 227488 346350 227808 346384
rect 227488 346294 227558 346350
rect 227614 346294 227682 346350
rect 227738 346294 227808 346350
rect 227488 346226 227808 346294
rect 227488 346170 227558 346226
rect 227614 346170 227682 346226
rect 227738 346170 227808 346226
rect 227488 346102 227808 346170
rect 227488 346046 227558 346102
rect 227614 346046 227682 346102
rect 227738 346046 227808 346102
rect 227488 345978 227808 346046
rect 227488 345922 227558 345978
rect 227614 345922 227682 345978
rect 227738 345922 227808 345978
rect 227488 345888 227808 345922
rect 258208 346350 258528 346384
rect 258208 346294 258278 346350
rect 258334 346294 258402 346350
rect 258458 346294 258528 346350
rect 258208 346226 258528 346294
rect 258208 346170 258278 346226
rect 258334 346170 258402 346226
rect 258458 346170 258528 346226
rect 258208 346102 258528 346170
rect 258208 346046 258278 346102
rect 258334 346046 258402 346102
rect 258458 346046 258528 346102
rect 258208 345978 258528 346046
rect 258208 345922 258278 345978
rect 258334 345922 258402 345978
rect 258458 345922 258528 345978
rect 258208 345888 258528 345922
rect 288928 346350 289248 346384
rect 288928 346294 288998 346350
rect 289054 346294 289122 346350
rect 289178 346294 289248 346350
rect 288928 346226 289248 346294
rect 288928 346170 288998 346226
rect 289054 346170 289122 346226
rect 289178 346170 289248 346226
rect 288928 346102 289248 346170
rect 288928 346046 288998 346102
rect 289054 346046 289122 346102
rect 289178 346046 289248 346102
rect 288928 345978 289248 346046
rect 288928 345922 288998 345978
rect 289054 345922 289122 345978
rect 289178 345922 289248 345978
rect 288928 345888 289248 345922
rect 319648 346350 319968 346384
rect 319648 346294 319718 346350
rect 319774 346294 319842 346350
rect 319898 346294 319968 346350
rect 319648 346226 319968 346294
rect 319648 346170 319718 346226
rect 319774 346170 319842 346226
rect 319898 346170 319968 346226
rect 319648 346102 319968 346170
rect 319648 346046 319718 346102
rect 319774 346046 319842 346102
rect 319898 346046 319968 346102
rect 319648 345978 319968 346046
rect 319648 345922 319718 345978
rect 319774 345922 319842 345978
rect 319898 345922 319968 345978
rect 319648 345888 319968 345922
rect 350368 346350 350688 346384
rect 350368 346294 350438 346350
rect 350494 346294 350562 346350
rect 350618 346294 350688 346350
rect 350368 346226 350688 346294
rect 350368 346170 350438 346226
rect 350494 346170 350562 346226
rect 350618 346170 350688 346226
rect 350368 346102 350688 346170
rect 350368 346046 350438 346102
rect 350494 346046 350562 346102
rect 350618 346046 350688 346102
rect 350368 345978 350688 346046
rect 350368 345922 350438 345978
rect 350494 345922 350562 345978
rect 350618 345922 350688 345978
rect 350368 345888 350688 345922
rect 381088 346350 381408 346384
rect 381088 346294 381158 346350
rect 381214 346294 381282 346350
rect 381338 346294 381408 346350
rect 381088 346226 381408 346294
rect 381088 346170 381158 346226
rect 381214 346170 381282 346226
rect 381338 346170 381408 346226
rect 381088 346102 381408 346170
rect 381088 346046 381158 346102
rect 381214 346046 381282 346102
rect 381338 346046 381408 346102
rect 381088 345978 381408 346046
rect 381088 345922 381158 345978
rect 381214 345922 381282 345978
rect 381338 345922 381408 345978
rect 381088 345888 381408 345922
rect 411808 346350 412128 346384
rect 411808 346294 411878 346350
rect 411934 346294 412002 346350
rect 412058 346294 412128 346350
rect 411808 346226 412128 346294
rect 411808 346170 411878 346226
rect 411934 346170 412002 346226
rect 412058 346170 412128 346226
rect 411808 346102 412128 346170
rect 411808 346046 411878 346102
rect 411934 346046 412002 346102
rect 412058 346046 412128 346102
rect 411808 345978 412128 346046
rect 411808 345922 411878 345978
rect 411934 345922 412002 345978
rect 412058 345922 412128 345978
rect 411808 345888 412128 345922
rect 442528 346350 442848 346384
rect 442528 346294 442598 346350
rect 442654 346294 442722 346350
rect 442778 346294 442848 346350
rect 442528 346226 442848 346294
rect 442528 346170 442598 346226
rect 442654 346170 442722 346226
rect 442778 346170 442848 346226
rect 442528 346102 442848 346170
rect 442528 346046 442598 346102
rect 442654 346046 442722 346102
rect 442778 346046 442848 346102
rect 442528 345978 442848 346046
rect 442528 345922 442598 345978
rect 442654 345922 442722 345978
rect 442778 345922 442848 345978
rect 442528 345888 442848 345922
rect 473248 346350 473568 346384
rect 473248 346294 473318 346350
rect 473374 346294 473442 346350
rect 473498 346294 473568 346350
rect 473248 346226 473568 346294
rect 473248 346170 473318 346226
rect 473374 346170 473442 346226
rect 473498 346170 473568 346226
rect 473248 346102 473568 346170
rect 473248 346046 473318 346102
rect 473374 346046 473442 346102
rect 473498 346046 473568 346102
rect 473248 345978 473568 346046
rect 473248 345922 473318 345978
rect 473374 345922 473442 345978
rect 473498 345922 473568 345978
rect 473248 345888 473568 345922
rect 503968 346350 504288 346384
rect 503968 346294 504038 346350
rect 504094 346294 504162 346350
rect 504218 346294 504288 346350
rect 503968 346226 504288 346294
rect 503968 346170 504038 346226
rect 504094 346170 504162 346226
rect 504218 346170 504288 346226
rect 503968 346102 504288 346170
rect 503968 346046 504038 346102
rect 504094 346046 504162 346102
rect 504218 346046 504288 346102
rect 503968 345978 504288 346046
rect 503968 345922 504038 345978
rect 504094 345922 504162 345978
rect 504218 345922 504288 345978
rect 503968 345888 504288 345922
rect 534688 346350 535008 346384
rect 534688 346294 534758 346350
rect 534814 346294 534882 346350
rect 534938 346294 535008 346350
rect 534688 346226 535008 346294
rect 534688 346170 534758 346226
rect 534814 346170 534882 346226
rect 534938 346170 535008 346226
rect 534688 346102 535008 346170
rect 534688 346046 534758 346102
rect 534814 346046 534882 346102
rect 534938 346046 535008 346102
rect 534688 345978 535008 346046
rect 534688 345922 534758 345978
rect 534814 345922 534882 345978
rect 534938 345922 535008 345978
rect 534688 345888 535008 345922
rect 565408 346350 565728 346384
rect 565408 346294 565478 346350
rect 565534 346294 565602 346350
rect 565658 346294 565728 346350
rect 565408 346226 565728 346294
rect 565408 346170 565478 346226
rect 565534 346170 565602 346226
rect 565658 346170 565728 346226
rect 565408 346102 565728 346170
rect 565408 346046 565478 346102
rect 565534 346046 565602 346102
rect 565658 346046 565728 346102
rect 565408 345978 565728 346046
rect 565408 345922 565478 345978
rect 565534 345922 565602 345978
rect 565658 345922 565728 345978
rect 565408 345888 565728 345922
rect 27808 334350 28128 334384
rect 27808 334294 27878 334350
rect 27934 334294 28002 334350
rect 28058 334294 28128 334350
rect 27808 334226 28128 334294
rect 27808 334170 27878 334226
rect 27934 334170 28002 334226
rect 28058 334170 28128 334226
rect 27808 334102 28128 334170
rect 27808 334046 27878 334102
rect 27934 334046 28002 334102
rect 28058 334046 28128 334102
rect 27808 333978 28128 334046
rect 27808 333922 27878 333978
rect 27934 333922 28002 333978
rect 28058 333922 28128 333978
rect 27808 333888 28128 333922
rect 58528 334350 58848 334384
rect 58528 334294 58598 334350
rect 58654 334294 58722 334350
rect 58778 334294 58848 334350
rect 58528 334226 58848 334294
rect 58528 334170 58598 334226
rect 58654 334170 58722 334226
rect 58778 334170 58848 334226
rect 58528 334102 58848 334170
rect 58528 334046 58598 334102
rect 58654 334046 58722 334102
rect 58778 334046 58848 334102
rect 58528 333978 58848 334046
rect 58528 333922 58598 333978
rect 58654 333922 58722 333978
rect 58778 333922 58848 333978
rect 58528 333888 58848 333922
rect 89248 334350 89568 334384
rect 89248 334294 89318 334350
rect 89374 334294 89442 334350
rect 89498 334294 89568 334350
rect 89248 334226 89568 334294
rect 89248 334170 89318 334226
rect 89374 334170 89442 334226
rect 89498 334170 89568 334226
rect 89248 334102 89568 334170
rect 89248 334046 89318 334102
rect 89374 334046 89442 334102
rect 89498 334046 89568 334102
rect 89248 333978 89568 334046
rect 89248 333922 89318 333978
rect 89374 333922 89442 333978
rect 89498 333922 89568 333978
rect 89248 333888 89568 333922
rect 119968 334350 120288 334384
rect 119968 334294 120038 334350
rect 120094 334294 120162 334350
rect 120218 334294 120288 334350
rect 119968 334226 120288 334294
rect 119968 334170 120038 334226
rect 120094 334170 120162 334226
rect 120218 334170 120288 334226
rect 119968 334102 120288 334170
rect 119968 334046 120038 334102
rect 120094 334046 120162 334102
rect 120218 334046 120288 334102
rect 119968 333978 120288 334046
rect 119968 333922 120038 333978
rect 120094 333922 120162 333978
rect 120218 333922 120288 333978
rect 119968 333888 120288 333922
rect 150688 334350 151008 334384
rect 150688 334294 150758 334350
rect 150814 334294 150882 334350
rect 150938 334294 151008 334350
rect 150688 334226 151008 334294
rect 150688 334170 150758 334226
rect 150814 334170 150882 334226
rect 150938 334170 151008 334226
rect 150688 334102 151008 334170
rect 150688 334046 150758 334102
rect 150814 334046 150882 334102
rect 150938 334046 151008 334102
rect 150688 333978 151008 334046
rect 150688 333922 150758 333978
rect 150814 333922 150882 333978
rect 150938 333922 151008 333978
rect 150688 333888 151008 333922
rect 181408 334350 181728 334384
rect 181408 334294 181478 334350
rect 181534 334294 181602 334350
rect 181658 334294 181728 334350
rect 181408 334226 181728 334294
rect 181408 334170 181478 334226
rect 181534 334170 181602 334226
rect 181658 334170 181728 334226
rect 181408 334102 181728 334170
rect 181408 334046 181478 334102
rect 181534 334046 181602 334102
rect 181658 334046 181728 334102
rect 181408 333978 181728 334046
rect 181408 333922 181478 333978
rect 181534 333922 181602 333978
rect 181658 333922 181728 333978
rect 181408 333888 181728 333922
rect 212128 334350 212448 334384
rect 212128 334294 212198 334350
rect 212254 334294 212322 334350
rect 212378 334294 212448 334350
rect 212128 334226 212448 334294
rect 212128 334170 212198 334226
rect 212254 334170 212322 334226
rect 212378 334170 212448 334226
rect 212128 334102 212448 334170
rect 212128 334046 212198 334102
rect 212254 334046 212322 334102
rect 212378 334046 212448 334102
rect 212128 333978 212448 334046
rect 212128 333922 212198 333978
rect 212254 333922 212322 333978
rect 212378 333922 212448 333978
rect 212128 333888 212448 333922
rect 242848 334350 243168 334384
rect 242848 334294 242918 334350
rect 242974 334294 243042 334350
rect 243098 334294 243168 334350
rect 242848 334226 243168 334294
rect 242848 334170 242918 334226
rect 242974 334170 243042 334226
rect 243098 334170 243168 334226
rect 242848 334102 243168 334170
rect 242848 334046 242918 334102
rect 242974 334046 243042 334102
rect 243098 334046 243168 334102
rect 242848 333978 243168 334046
rect 242848 333922 242918 333978
rect 242974 333922 243042 333978
rect 243098 333922 243168 333978
rect 242848 333888 243168 333922
rect 273568 334350 273888 334384
rect 273568 334294 273638 334350
rect 273694 334294 273762 334350
rect 273818 334294 273888 334350
rect 273568 334226 273888 334294
rect 273568 334170 273638 334226
rect 273694 334170 273762 334226
rect 273818 334170 273888 334226
rect 273568 334102 273888 334170
rect 273568 334046 273638 334102
rect 273694 334046 273762 334102
rect 273818 334046 273888 334102
rect 273568 333978 273888 334046
rect 273568 333922 273638 333978
rect 273694 333922 273762 333978
rect 273818 333922 273888 333978
rect 273568 333888 273888 333922
rect 304288 334350 304608 334384
rect 304288 334294 304358 334350
rect 304414 334294 304482 334350
rect 304538 334294 304608 334350
rect 304288 334226 304608 334294
rect 304288 334170 304358 334226
rect 304414 334170 304482 334226
rect 304538 334170 304608 334226
rect 304288 334102 304608 334170
rect 304288 334046 304358 334102
rect 304414 334046 304482 334102
rect 304538 334046 304608 334102
rect 304288 333978 304608 334046
rect 304288 333922 304358 333978
rect 304414 333922 304482 333978
rect 304538 333922 304608 333978
rect 304288 333888 304608 333922
rect 335008 334350 335328 334384
rect 335008 334294 335078 334350
rect 335134 334294 335202 334350
rect 335258 334294 335328 334350
rect 335008 334226 335328 334294
rect 335008 334170 335078 334226
rect 335134 334170 335202 334226
rect 335258 334170 335328 334226
rect 335008 334102 335328 334170
rect 335008 334046 335078 334102
rect 335134 334046 335202 334102
rect 335258 334046 335328 334102
rect 335008 333978 335328 334046
rect 335008 333922 335078 333978
rect 335134 333922 335202 333978
rect 335258 333922 335328 333978
rect 335008 333888 335328 333922
rect 365728 334350 366048 334384
rect 365728 334294 365798 334350
rect 365854 334294 365922 334350
rect 365978 334294 366048 334350
rect 365728 334226 366048 334294
rect 365728 334170 365798 334226
rect 365854 334170 365922 334226
rect 365978 334170 366048 334226
rect 365728 334102 366048 334170
rect 365728 334046 365798 334102
rect 365854 334046 365922 334102
rect 365978 334046 366048 334102
rect 365728 333978 366048 334046
rect 365728 333922 365798 333978
rect 365854 333922 365922 333978
rect 365978 333922 366048 333978
rect 365728 333888 366048 333922
rect 396448 334350 396768 334384
rect 396448 334294 396518 334350
rect 396574 334294 396642 334350
rect 396698 334294 396768 334350
rect 396448 334226 396768 334294
rect 396448 334170 396518 334226
rect 396574 334170 396642 334226
rect 396698 334170 396768 334226
rect 396448 334102 396768 334170
rect 396448 334046 396518 334102
rect 396574 334046 396642 334102
rect 396698 334046 396768 334102
rect 396448 333978 396768 334046
rect 396448 333922 396518 333978
rect 396574 333922 396642 333978
rect 396698 333922 396768 333978
rect 396448 333888 396768 333922
rect 427168 334350 427488 334384
rect 427168 334294 427238 334350
rect 427294 334294 427362 334350
rect 427418 334294 427488 334350
rect 427168 334226 427488 334294
rect 427168 334170 427238 334226
rect 427294 334170 427362 334226
rect 427418 334170 427488 334226
rect 427168 334102 427488 334170
rect 427168 334046 427238 334102
rect 427294 334046 427362 334102
rect 427418 334046 427488 334102
rect 427168 333978 427488 334046
rect 427168 333922 427238 333978
rect 427294 333922 427362 333978
rect 427418 333922 427488 333978
rect 427168 333888 427488 333922
rect 457888 334350 458208 334384
rect 457888 334294 457958 334350
rect 458014 334294 458082 334350
rect 458138 334294 458208 334350
rect 457888 334226 458208 334294
rect 457888 334170 457958 334226
rect 458014 334170 458082 334226
rect 458138 334170 458208 334226
rect 457888 334102 458208 334170
rect 457888 334046 457958 334102
rect 458014 334046 458082 334102
rect 458138 334046 458208 334102
rect 457888 333978 458208 334046
rect 457888 333922 457958 333978
rect 458014 333922 458082 333978
rect 458138 333922 458208 333978
rect 457888 333888 458208 333922
rect 488608 334350 488928 334384
rect 488608 334294 488678 334350
rect 488734 334294 488802 334350
rect 488858 334294 488928 334350
rect 488608 334226 488928 334294
rect 488608 334170 488678 334226
rect 488734 334170 488802 334226
rect 488858 334170 488928 334226
rect 488608 334102 488928 334170
rect 488608 334046 488678 334102
rect 488734 334046 488802 334102
rect 488858 334046 488928 334102
rect 488608 333978 488928 334046
rect 488608 333922 488678 333978
rect 488734 333922 488802 333978
rect 488858 333922 488928 333978
rect 488608 333888 488928 333922
rect 519328 334350 519648 334384
rect 519328 334294 519398 334350
rect 519454 334294 519522 334350
rect 519578 334294 519648 334350
rect 519328 334226 519648 334294
rect 519328 334170 519398 334226
rect 519454 334170 519522 334226
rect 519578 334170 519648 334226
rect 519328 334102 519648 334170
rect 519328 334046 519398 334102
rect 519454 334046 519522 334102
rect 519578 334046 519648 334102
rect 519328 333978 519648 334046
rect 519328 333922 519398 333978
rect 519454 333922 519522 333978
rect 519578 333922 519648 333978
rect 519328 333888 519648 333922
rect 550048 334350 550368 334384
rect 550048 334294 550118 334350
rect 550174 334294 550242 334350
rect 550298 334294 550368 334350
rect 550048 334226 550368 334294
rect 550048 334170 550118 334226
rect 550174 334170 550242 334226
rect 550298 334170 550368 334226
rect 550048 334102 550368 334170
rect 550048 334046 550118 334102
rect 550174 334046 550242 334102
rect 550298 334046 550368 334102
rect 550048 333978 550368 334046
rect 550048 333922 550118 333978
rect 550174 333922 550242 333978
rect 550298 333922 550368 333978
rect 550048 333888 550368 333922
rect 6188 333442 6244 333452
rect 5418 328294 5514 328350
rect 5570 328294 5638 328350
rect 5694 328294 5762 328350
rect 5818 328294 5886 328350
rect 5942 328294 6038 328350
rect 5418 328226 6038 328294
rect 5418 328170 5514 328226
rect 5570 328170 5638 328226
rect 5694 328170 5762 328226
rect 5818 328170 5886 328226
rect 5942 328170 6038 328226
rect 5418 328102 6038 328170
rect 5418 328046 5514 328102
rect 5570 328046 5638 328102
rect 5694 328046 5762 328102
rect 5818 328046 5886 328102
rect 5942 328046 6038 328102
rect 5418 327978 6038 328046
rect 5418 327922 5514 327978
rect 5570 327922 5638 327978
rect 5694 327922 5762 327978
rect 5818 327922 5886 327978
rect 5942 327922 6038 327978
rect 4172 312386 4228 312396
rect 4284 319060 4340 319070
rect -956 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 -336 310350
rect -956 310226 -336 310294
rect -956 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 -336 310226
rect -956 310102 -336 310170
rect -956 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 -336 310102
rect -956 309978 -336 310046
rect -956 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 -336 309978
rect -956 292350 -336 309922
rect 4284 301924 4340 319004
rect 4284 301858 4340 301868
rect 5418 310350 6038 327922
rect 12448 328350 12768 328384
rect 12448 328294 12518 328350
rect 12574 328294 12642 328350
rect 12698 328294 12768 328350
rect 12448 328226 12768 328294
rect 12448 328170 12518 328226
rect 12574 328170 12642 328226
rect 12698 328170 12768 328226
rect 12448 328102 12768 328170
rect 12448 328046 12518 328102
rect 12574 328046 12642 328102
rect 12698 328046 12768 328102
rect 12448 327978 12768 328046
rect 12448 327922 12518 327978
rect 12574 327922 12642 327978
rect 12698 327922 12768 327978
rect 12448 327888 12768 327922
rect 43168 328350 43488 328384
rect 43168 328294 43238 328350
rect 43294 328294 43362 328350
rect 43418 328294 43488 328350
rect 43168 328226 43488 328294
rect 43168 328170 43238 328226
rect 43294 328170 43362 328226
rect 43418 328170 43488 328226
rect 43168 328102 43488 328170
rect 43168 328046 43238 328102
rect 43294 328046 43362 328102
rect 43418 328046 43488 328102
rect 43168 327978 43488 328046
rect 43168 327922 43238 327978
rect 43294 327922 43362 327978
rect 43418 327922 43488 327978
rect 43168 327888 43488 327922
rect 73888 328350 74208 328384
rect 73888 328294 73958 328350
rect 74014 328294 74082 328350
rect 74138 328294 74208 328350
rect 73888 328226 74208 328294
rect 73888 328170 73958 328226
rect 74014 328170 74082 328226
rect 74138 328170 74208 328226
rect 73888 328102 74208 328170
rect 73888 328046 73958 328102
rect 74014 328046 74082 328102
rect 74138 328046 74208 328102
rect 73888 327978 74208 328046
rect 73888 327922 73958 327978
rect 74014 327922 74082 327978
rect 74138 327922 74208 327978
rect 73888 327888 74208 327922
rect 104608 328350 104928 328384
rect 104608 328294 104678 328350
rect 104734 328294 104802 328350
rect 104858 328294 104928 328350
rect 104608 328226 104928 328294
rect 104608 328170 104678 328226
rect 104734 328170 104802 328226
rect 104858 328170 104928 328226
rect 104608 328102 104928 328170
rect 104608 328046 104678 328102
rect 104734 328046 104802 328102
rect 104858 328046 104928 328102
rect 104608 327978 104928 328046
rect 104608 327922 104678 327978
rect 104734 327922 104802 327978
rect 104858 327922 104928 327978
rect 104608 327888 104928 327922
rect 135328 328350 135648 328384
rect 135328 328294 135398 328350
rect 135454 328294 135522 328350
rect 135578 328294 135648 328350
rect 135328 328226 135648 328294
rect 135328 328170 135398 328226
rect 135454 328170 135522 328226
rect 135578 328170 135648 328226
rect 135328 328102 135648 328170
rect 135328 328046 135398 328102
rect 135454 328046 135522 328102
rect 135578 328046 135648 328102
rect 135328 327978 135648 328046
rect 135328 327922 135398 327978
rect 135454 327922 135522 327978
rect 135578 327922 135648 327978
rect 135328 327888 135648 327922
rect 166048 328350 166368 328384
rect 166048 328294 166118 328350
rect 166174 328294 166242 328350
rect 166298 328294 166368 328350
rect 166048 328226 166368 328294
rect 166048 328170 166118 328226
rect 166174 328170 166242 328226
rect 166298 328170 166368 328226
rect 166048 328102 166368 328170
rect 166048 328046 166118 328102
rect 166174 328046 166242 328102
rect 166298 328046 166368 328102
rect 166048 327978 166368 328046
rect 166048 327922 166118 327978
rect 166174 327922 166242 327978
rect 166298 327922 166368 327978
rect 166048 327888 166368 327922
rect 196768 328350 197088 328384
rect 196768 328294 196838 328350
rect 196894 328294 196962 328350
rect 197018 328294 197088 328350
rect 196768 328226 197088 328294
rect 196768 328170 196838 328226
rect 196894 328170 196962 328226
rect 197018 328170 197088 328226
rect 196768 328102 197088 328170
rect 196768 328046 196838 328102
rect 196894 328046 196962 328102
rect 197018 328046 197088 328102
rect 196768 327978 197088 328046
rect 196768 327922 196838 327978
rect 196894 327922 196962 327978
rect 197018 327922 197088 327978
rect 196768 327888 197088 327922
rect 227488 328350 227808 328384
rect 227488 328294 227558 328350
rect 227614 328294 227682 328350
rect 227738 328294 227808 328350
rect 227488 328226 227808 328294
rect 227488 328170 227558 328226
rect 227614 328170 227682 328226
rect 227738 328170 227808 328226
rect 227488 328102 227808 328170
rect 227488 328046 227558 328102
rect 227614 328046 227682 328102
rect 227738 328046 227808 328102
rect 227488 327978 227808 328046
rect 227488 327922 227558 327978
rect 227614 327922 227682 327978
rect 227738 327922 227808 327978
rect 227488 327888 227808 327922
rect 258208 328350 258528 328384
rect 258208 328294 258278 328350
rect 258334 328294 258402 328350
rect 258458 328294 258528 328350
rect 258208 328226 258528 328294
rect 258208 328170 258278 328226
rect 258334 328170 258402 328226
rect 258458 328170 258528 328226
rect 258208 328102 258528 328170
rect 258208 328046 258278 328102
rect 258334 328046 258402 328102
rect 258458 328046 258528 328102
rect 258208 327978 258528 328046
rect 258208 327922 258278 327978
rect 258334 327922 258402 327978
rect 258458 327922 258528 327978
rect 258208 327888 258528 327922
rect 288928 328350 289248 328384
rect 288928 328294 288998 328350
rect 289054 328294 289122 328350
rect 289178 328294 289248 328350
rect 288928 328226 289248 328294
rect 288928 328170 288998 328226
rect 289054 328170 289122 328226
rect 289178 328170 289248 328226
rect 288928 328102 289248 328170
rect 288928 328046 288998 328102
rect 289054 328046 289122 328102
rect 289178 328046 289248 328102
rect 288928 327978 289248 328046
rect 288928 327922 288998 327978
rect 289054 327922 289122 327978
rect 289178 327922 289248 327978
rect 288928 327888 289248 327922
rect 319648 328350 319968 328384
rect 319648 328294 319718 328350
rect 319774 328294 319842 328350
rect 319898 328294 319968 328350
rect 319648 328226 319968 328294
rect 319648 328170 319718 328226
rect 319774 328170 319842 328226
rect 319898 328170 319968 328226
rect 319648 328102 319968 328170
rect 319648 328046 319718 328102
rect 319774 328046 319842 328102
rect 319898 328046 319968 328102
rect 319648 327978 319968 328046
rect 319648 327922 319718 327978
rect 319774 327922 319842 327978
rect 319898 327922 319968 327978
rect 319648 327888 319968 327922
rect 350368 328350 350688 328384
rect 350368 328294 350438 328350
rect 350494 328294 350562 328350
rect 350618 328294 350688 328350
rect 350368 328226 350688 328294
rect 350368 328170 350438 328226
rect 350494 328170 350562 328226
rect 350618 328170 350688 328226
rect 350368 328102 350688 328170
rect 350368 328046 350438 328102
rect 350494 328046 350562 328102
rect 350618 328046 350688 328102
rect 350368 327978 350688 328046
rect 350368 327922 350438 327978
rect 350494 327922 350562 327978
rect 350618 327922 350688 327978
rect 350368 327888 350688 327922
rect 381088 328350 381408 328384
rect 381088 328294 381158 328350
rect 381214 328294 381282 328350
rect 381338 328294 381408 328350
rect 381088 328226 381408 328294
rect 381088 328170 381158 328226
rect 381214 328170 381282 328226
rect 381338 328170 381408 328226
rect 381088 328102 381408 328170
rect 381088 328046 381158 328102
rect 381214 328046 381282 328102
rect 381338 328046 381408 328102
rect 381088 327978 381408 328046
rect 381088 327922 381158 327978
rect 381214 327922 381282 327978
rect 381338 327922 381408 327978
rect 381088 327888 381408 327922
rect 411808 328350 412128 328384
rect 411808 328294 411878 328350
rect 411934 328294 412002 328350
rect 412058 328294 412128 328350
rect 411808 328226 412128 328294
rect 411808 328170 411878 328226
rect 411934 328170 412002 328226
rect 412058 328170 412128 328226
rect 411808 328102 412128 328170
rect 411808 328046 411878 328102
rect 411934 328046 412002 328102
rect 412058 328046 412128 328102
rect 411808 327978 412128 328046
rect 411808 327922 411878 327978
rect 411934 327922 412002 327978
rect 412058 327922 412128 327978
rect 411808 327888 412128 327922
rect 442528 328350 442848 328384
rect 442528 328294 442598 328350
rect 442654 328294 442722 328350
rect 442778 328294 442848 328350
rect 442528 328226 442848 328294
rect 442528 328170 442598 328226
rect 442654 328170 442722 328226
rect 442778 328170 442848 328226
rect 442528 328102 442848 328170
rect 442528 328046 442598 328102
rect 442654 328046 442722 328102
rect 442778 328046 442848 328102
rect 442528 327978 442848 328046
rect 442528 327922 442598 327978
rect 442654 327922 442722 327978
rect 442778 327922 442848 327978
rect 442528 327888 442848 327922
rect 473248 328350 473568 328384
rect 473248 328294 473318 328350
rect 473374 328294 473442 328350
rect 473498 328294 473568 328350
rect 473248 328226 473568 328294
rect 473248 328170 473318 328226
rect 473374 328170 473442 328226
rect 473498 328170 473568 328226
rect 473248 328102 473568 328170
rect 473248 328046 473318 328102
rect 473374 328046 473442 328102
rect 473498 328046 473568 328102
rect 473248 327978 473568 328046
rect 473248 327922 473318 327978
rect 473374 327922 473442 327978
rect 473498 327922 473568 327978
rect 473248 327888 473568 327922
rect 503968 328350 504288 328384
rect 503968 328294 504038 328350
rect 504094 328294 504162 328350
rect 504218 328294 504288 328350
rect 503968 328226 504288 328294
rect 503968 328170 504038 328226
rect 504094 328170 504162 328226
rect 504218 328170 504288 328226
rect 503968 328102 504288 328170
rect 503968 328046 504038 328102
rect 504094 328046 504162 328102
rect 504218 328046 504288 328102
rect 503968 327978 504288 328046
rect 503968 327922 504038 327978
rect 504094 327922 504162 327978
rect 504218 327922 504288 327978
rect 503968 327888 504288 327922
rect 534688 328350 535008 328384
rect 534688 328294 534758 328350
rect 534814 328294 534882 328350
rect 534938 328294 535008 328350
rect 534688 328226 535008 328294
rect 534688 328170 534758 328226
rect 534814 328170 534882 328226
rect 534938 328170 535008 328226
rect 534688 328102 535008 328170
rect 534688 328046 534758 328102
rect 534814 328046 534882 328102
rect 534938 328046 535008 328102
rect 534688 327978 535008 328046
rect 534688 327922 534758 327978
rect 534814 327922 534882 327978
rect 534938 327922 535008 327978
rect 534688 327888 535008 327922
rect 565408 328350 565728 328384
rect 565408 328294 565478 328350
rect 565534 328294 565602 328350
rect 565658 328294 565728 328350
rect 565408 328226 565728 328294
rect 565408 328170 565478 328226
rect 565534 328170 565602 328226
rect 565658 328170 565728 328226
rect 565408 328102 565728 328170
rect 565408 328046 565478 328102
rect 565534 328046 565602 328102
rect 565658 328046 565728 328102
rect 565408 327978 565728 328046
rect 565408 327922 565478 327978
rect 565534 327922 565602 327978
rect 565658 327922 565728 327978
rect 565408 327888 565728 327922
rect 585452 318276 585508 350700
rect 585676 350532 585732 377132
rect 585676 350466 585732 350476
rect 589098 364350 589718 381922
rect 589098 364294 589194 364350
rect 589250 364294 589318 364350
rect 589374 364294 589442 364350
rect 589498 364294 589566 364350
rect 589622 364294 589718 364350
rect 589098 364226 589718 364294
rect 589098 364170 589194 364226
rect 589250 364170 589318 364226
rect 589374 364170 589442 364226
rect 589498 364170 589566 364226
rect 589622 364170 589718 364226
rect 589098 364102 589718 364170
rect 589098 364046 589194 364102
rect 589250 364046 589318 364102
rect 589374 364046 589442 364102
rect 589498 364046 589566 364102
rect 589622 364046 589718 364102
rect 589098 363978 589718 364046
rect 592818 424350 593438 441922
rect 592818 424294 592914 424350
rect 592970 424294 593038 424350
rect 593094 424294 593162 424350
rect 593218 424294 593286 424350
rect 593342 424294 593438 424350
rect 592818 424226 593438 424294
rect 592818 424170 592914 424226
rect 592970 424170 593038 424226
rect 593094 424170 593162 424226
rect 593218 424170 593286 424226
rect 593342 424170 593438 424226
rect 592818 424102 593438 424170
rect 592818 424046 592914 424102
rect 592970 424046 593038 424102
rect 593094 424046 593162 424102
rect 593218 424046 593286 424102
rect 593342 424046 593438 424102
rect 592818 423978 593438 424046
rect 592818 423922 592914 423978
rect 592970 423922 593038 423978
rect 593094 423922 593162 423978
rect 593218 423922 593286 423978
rect 593342 423922 593438 423978
rect 592818 406350 593438 423922
rect 592818 406294 592914 406350
rect 592970 406294 593038 406350
rect 593094 406294 593162 406350
rect 593218 406294 593286 406350
rect 593342 406294 593438 406350
rect 592818 406226 593438 406294
rect 592818 406170 592914 406226
rect 592970 406170 593038 406226
rect 593094 406170 593162 406226
rect 593218 406170 593286 406226
rect 593342 406170 593438 406226
rect 592818 406102 593438 406170
rect 592818 406046 592914 406102
rect 592970 406046 593038 406102
rect 593094 406046 593162 406102
rect 593218 406046 593286 406102
rect 593342 406046 593438 406102
rect 592818 405978 593438 406046
rect 592818 405922 592914 405978
rect 592970 405922 593038 405978
rect 593094 405922 593162 405978
rect 593218 405922 593286 405978
rect 593342 405922 593438 405978
rect 592818 388350 593438 405922
rect 592818 388294 592914 388350
rect 592970 388294 593038 388350
rect 593094 388294 593162 388350
rect 593218 388294 593286 388350
rect 593342 388294 593438 388350
rect 592818 388226 593438 388294
rect 592818 388170 592914 388226
rect 592970 388170 593038 388226
rect 593094 388170 593162 388226
rect 593218 388170 593286 388226
rect 593342 388170 593438 388226
rect 592818 388102 593438 388170
rect 592818 388046 592914 388102
rect 592970 388046 593038 388102
rect 593094 388046 593162 388102
rect 593218 388046 593286 388102
rect 593342 388046 593438 388102
rect 592818 387978 593438 388046
rect 592818 387922 592914 387978
rect 592970 387922 593038 387978
rect 593094 387922 593162 387978
rect 593218 387922 593286 387978
rect 593342 387922 593438 387978
rect 592818 370350 593438 387922
rect 592818 370294 592914 370350
rect 592970 370294 593038 370350
rect 593094 370294 593162 370350
rect 593218 370294 593286 370350
rect 593342 370294 593438 370350
rect 592818 370226 593438 370294
rect 592818 370170 592914 370226
rect 592970 370170 593038 370226
rect 593094 370170 593162 370226
rect 593218 370170 593286 370226
rect 593342 370170 593438 370226
rect 592818 370102 593438 370170
rect 592818 370046 592914 370102
rect 592970 370046 593038 370102
rect 593094 370046 593162 370102
rect 593218 370046 593286 370102
rect 593342 370046 593438 370102
rect 592818 369978 593438 370046
rect 592818 369922 592914 369978
rect 592970 369922 593038 369978
rect 593094 369922 593162 369978
rect 593218 369922 593286 369978
rect 593342 369922 593438 369978
rect 589098 363922 589194 363978
rect 589250 363922 589318 363978
rect 589374 363922 589442 363978
rect 589498 363922 589566 363978
rect 589622 363922 589718 363978
rect 589098 346350 589718 363922
rect 589098 346294 589194 346350
rect 589250 346294 589318 346350
rect 589374 346294 589442 346350
rect 589498 346294 589566 346350
rect 589622 346294 589718 346350
rect 589098 346226 589718 346294
rect 589098 346170 589194 346226
rect 589250 346170 589318 346226
rect 589374 346170 589442 346226
rect 589498 346170 589566 346226
rect 589622 346170 589718 346226
rect 589098 346102 589718 346170
rect 589098 346046 589194 346102
rect 589250 346046 589318 346102
rect 589374 346046 589442 346102
rect 589498 346046 589566 346102
rect 589622 346046 589718 346102
rect 589098 345978 589718 346046
rect 589098 345922 589194 345978
rect 589250 345922 589318 345978
rect 589374 345922 589442 345978
rect 589498 345922 589566 345978
rect 589622 345922 589718 345978
rect 585676 337540 585732 337550
rect 585452 318210 585508 318220
rect 585564 324324 585620 324334
rect 27808 316350 28128 316384
rect 27808 316294 27878 316350
rect 27934 316294 28002 316350
rect 28058 316294 28128 316350
rect 27808 316226 28128 316294
rect 27808 316170 27878 316226
rect 27934 316170 28002 316226
rect 28058 316170 28128 316226
rect 27808 316102 28128 316170
rect 27808 316046 27878 316102
rect 27934 316046 28002 316102
rect 28058 316046 28128 316102
rect 27808 315978 28128 316046
rect 27808 315922 27878 315978
rect 27934 315922 28002 315978
rect 28058 315922 28128 315978
rect 27808 315888 28128 315922
rect 58528 316350 58848 316384
rect 58528 316294 58598 316350
rect 58654 316294 58722 316350
rect 58778 316294 58848 316350
rect 58528 316226 58848 316294
rect 58528 316170 58598 316226
rect 58654 316170 58722 316226
rect 58778 316170 58848 316226
rect 58528 316102 58848 316170
rect 58528 316046 58598 316102
rect 58654 316046 58722 316102
rect 58778 316046 58848 316102
rect 58528 315978 58848 316046
rect 58528 315922 58598 315978
rect 58654 315922 58722 315978
rect 58778 315922 58848 315978
rect 58528 315888 58848 315922
rect 89248 316350 89568 316384
rect 89248 316294 89318 316350
rect 89374 316294 89442 316350
rect 89498 316294 89568 316350
rect 89248 316226 89568 316294
rect 89248 316170 89318 316226
rect 89374 316170 89442 316226
rect 89498 316170 89568 316226
rect 89248 316102 89568 316170
rect 89248 316046 89318 316102
rect 89374 316046 89442 316102
rect 89498 316046 89568 316102
rect 89248 315978 89568 316046
rect 89248 315922 89318 315978
rect 89374 315922 89442 315978
rect 89498 315922 89568 315978
rect 89248 315888 89568 315922
rect 119968 316350 120288 316384
rect 119968 316294 120038 316350
rect 120094 316294 120162 316350
rect 120218 316294 120288 316350
rect 119968 316226 120288 316294
rect 119968 316170 120038 316226
rect 120094 316170 120162 316226
rect 120218 316170 120288 316226
rect 119968 316102 120288 316170
rect 119968 316046 120038 316102
rect 120094 316046 120162 316102
rect 120218 316046 120288 316102
rect 119968 315978 120288 316046
rect 119968 315922 120038 315978
rect 120094 315922 120162 315978
rect 120218 315922 120288 315978
rect 119968 315888 120288 315922
rect 150688 316350 151008 316384
rect 150688 316294 150758 316350
rect 150814 316294 150882 316350
rect 150938 316294 151008 316350
rect 150688 316226 151008 316294
rect 150688 316170 150758 316226
rect 150814 316170 150882 316226
rect 150938 316170 151008 316226
rect 150688 316102 151008 316170
rect 150688 316046 150758 316102
rect 150814 316046 150882 316102
rect 150938 316046 151008 316102
rect 150688 315978 151008 316046
rect 150688 315922 150758 315978
rect 150814 315922 150882 315978
rect 150938 315922 151008 315978
rect 150688 315888 151008 315922
rect 181408 316350 181728 316384
rect 181408 316294 181478 316350
rect 181534 316294 181602 316350
rect 181658 316294 181728 316350
rect 181408 316226 181728 316294
rect 181408 316170 181478 316226
rect 181534 316170 181602 316226
rect 181658 316170 181728 316226
rect 181408 316102 181728 316170
rect 181408 316046 181478 316102
rect 181534 316046 181602 316102
rect 181658 316046 181728 316102
rect 181408 315978 181728 316046
rect 181408 315922 181478 315978
rect 181534 315922 181602 315978
rect 181658 315922 181728 315978
rect 181408 315888 181728 315922
rect 212128 316350 212448 316384
rect 212128 316294 212198 316350
rect 212254 316294 212322 316350
rect 212378 316294 212448 316350
rect 212128 316226 212448 316294
rect 212128 316170 212198 316226
rect 212254 316170 212322 316226
rect 212378 316170 212448 316226
rect 212128 316102 212448 316170
rect 212128 316046 212198 316102
rect 212254 316046 212322 316102
rect 212378 316046 212448 316102
rect 212128 315978 212448 316046
rect 212128 315922 212198 315978
rect 212254 315922 212322 315978
rect 212378 315922 212448 315978
rect 212128 315888 212448 315922
rect 242848 316350 243168 316384
rect 242848 316294 242918 316350
rect 242974 316294 243042 316350
rect 243098 316294 243168 316350
rect 242848 316226 243168 316294
rect 242848 316170 242918 316226
rect 242974 316170 243042 316226
rect 243098 316170 243168 316226
rect 242848 316102 243168 316170
rect 242848 316046 242918 316102
rect 242974 316046 243042 316102
rect 243098 316046 243168 316102
rect 242848 315978 243168 316046
rect 242848 315922 242918 315978
rect 242974 315922 243042 315978
rect 243098 315922 243168 315978
rect 242848 315888 243168 315922
rect 273568 316350 273888 316384
rect 273568 316294 273638 316350
rect 273694 316294 273762 316350
rect 273818 316294 273888 316350
rect 273568 316226 273888 316294
rect 273568 316170 273638 316226
rect 273694 316170 273762 316226
rect 273818 316170 273888 316226
rect 273568 316102 273888 316170
rect 273568 316046 273638 316102
rect 273694 316046 273762 316102
rect 273818 316046 273888 316102
rect 273568 315978 273888 316046
rect 273568 315922 273638 315978
rect 273694 315922 273762 315978
rect 273818 315922 273888 315978
rect 273568 315888 273888 315922
rect 304288 316350 304608 316384
rect 304288 316294 304358 316350
rect 304414 316294 304482 316350
rect 304538 316294 304608 316350
rect 304288 316226 304608 316294
rect 304288 316170 304358 316226
rect 304414 316170 304482 316226
rect 304538 316170 304608 316226
rect 304288 316102 304608 316170
rect 304288 316046 304358 316102
rect 304414 316046 304482 316102
rect 304538 316046 304608 316102
rect 304288 315978 304608 316046
rect 304288 315922 304358 315978
rect 304414 315922 304482 315978
rect 304538 315922 304608 315978
rect 304288 315888 304608 315922
rect 335008 316350 335328 316384
rect 335008 316294 335078 316350
rect 335134 316294 335202 316350
rect 335258 316294 335328 316350
rect 335008 316226 335328 316294
rect 335008 316170 335078 316226
rect 335134 316170 335202 316226
rect 335258 316170 335328 316226
rect 335008 316102 335328 316170
rect 335008 316046 335078 316102
rect 335134 316046 335202 316102
rect 335258 316046 335328 316102
rect 335008 315978 335328 316046
rect 335008 315922 335078 315978
rect 335134 315922 335202 315978
rect 335258 315922 335328 315978
rect 335008 315888 335328 315922
rect 365728 316350 366048 316384
rect 365728 316294 365798 316350
rect 365854 316294 365922 316350
rect 365978 316294 366048 316350
rect 365728 316226 366048 316294
rect 365728 316170 365798 316226
rect 365854 316170 365922 316226
rect 365978 316170 366048 316226
rect 365728 316102 366048 316170
rect 365728 316046 365798 316102
rect 365854 316046 365922 316102
rect 365978 316046 366048 316102
rect 365728 315978 366048 316046
rect 365728 315922 365798 315978
rect 365854 315922 365922 315978
rect 365978 315922 366048 315978
rect 365728 315888 366048 315922
rect 396448 316350 396768 316384
rect 396448 316294 396518 316350
rect 396574 316294 396642 316350
rect 396698 316294 396768 316350
rect 396448 316226 396768 316294
rect 396448 316170 396518 316226
rect 396574 316170 396642 316226
rect 396698 316170 396768 316226
rect 396448 316102 396768 316170
rect 396448 316046 396518 316102
rect 396574 316046 396642 316102
rect 396698 316046 396768 316102
rect 396448 315978 396768 316046
rect 396448 315922 396518 315978
rect 396574 315922 396642 315978
rect 396698 315922 396768 315978
rect 396448 315888 396768 315922
rect 427168 316350 427488 316384
rect 427168 316294 427238 316350
rect 427294 316294 427362 316350
rect 427418 316294 427488 316350
rect 427168 316226 427488 316294
rect 427168 316170 427238 316226
rect 427294 316170 427362 316226
rect 427418 316170 427488 316226
rect 427168 316102 427488 316170
rect 427168 316046 427238 316102
rect 427294 316046 427362 316102
rect 427418 316046 427488 316102
rect 427168 315978 427488 316046
rect 427168 315922 427238 315978
rect 427294 315922 427362 315978
rect 427418 315922 427488 315978
rect 427168 315888 427488 315922
rect 457888 316350 458208 316384
rect 457888 316294 457958 316350
rect 458014 316294 458082 316350
rect 458138 316294 458208 316350
rect 457888 316226 458208 316294
rect 457888 316170 457958 316226
rect 458014 316170 458082 316226
rect 458138 316170 458208 316226
rect 457888 316102 458208 316170
rect 457888 316046 457958 316102
rect 458014 316046 458082 316102
rect 458138 316046 458208 316102
rect 457888 315978 458208 316046
rect 457888 315922 457958 315978
rect 458014 315922 458082 315978
rect 458138 315922 458208 315978
rect 457888 315888 458208 315922
rect 488608 316350 488928 316384
rect 488608 316294 488678 316350
rect 488734 316294 488802 316350
rect 488858 316294 488928 316350
rect 488608 316226 488928 316294
rect 488608 316170 488678 316226
rect 488734 316170 488802 316226
rect 488858 316170 488928 316226
rect 488608 316102 488928 316170
rect 488608 316046 488678 316102
rect 488734 316046 488802 316102
rect 488858 316046 488928 316102
rect 488608 315978 488928 316046
rect 488608 315922 488678 315978
rect 488734 315922 488802 315978
rect 488858 315922 488928 315978
rect 488608 315888 488928 315922
rect 519328 316350 519648 316384
rect 519328 316294 519398 316350
rect 519454 316294 519522 316350
rect 519578 316294 519648 316350
rect 519328 316226 519648 316294
rect 519328 316170 519398 316226
rect 519454 316170 519522 316226
rect 519578 316170 519648 316226
rect 519328 316102 519648 316170
rect 519328 316046 519398 316102
rect 519454 316046 519522 316102
rect 519578 316046 519648 316102
rect 519328 315978 519648 316046
rect 519328 315922 519398 315978
rect 519454 315922 519522 315978
rect 519578 315922 519648 315978
rect 519328 315888 519648 315922
rect 550048 316350 550368 316384
rect 550048 316294 550118 316350
rect 550174 316294 550242 316350
rect 550298 316294 550368 316350
rect 550048 316226 550368 316294
rect 550048 316170 550118 316226
rect 550174 316170 550242 316226
rect 550298 316170 550368 316226
rect 550048 316102 550368 316170
rect 550048 316046 550118 316102
rect 550174 316046 550242 316102
rect 550298 316046 550368 316102
rect 550048 315978 550368 316046
rect 550048 315922 550118 315978
rect 550174 315922 550242 315978
rect 550298 315922 550368 315978
rect 550048 315888 550368 315922
rect 585452 311108 585508 311118
rect 5418 310294 5514 310350
rect 5570 310294 5638 310350
rect 5694 310294 5762 310350
rect 5818 310294 5886 310350
rect 5942 310294 6038 310350
rect 5418 310226 6038 310294
rect 5418 310170 5514 310226
rect 5570 310170 5638 310226
rect 5694 310170 5762 310226
rect 5818 310170 5886 310226
rect 5942 310170 6038 310226
rect 5418 310102 6038 310170
rect 5418 310046 5514 310102
rect 5570 310046 5638 310102
rect 5694 310046 5762 310102
rect 5818 310046 5886 310102
rect 5942 310046 6038 310102
rect 5418 309978 6038 310046
rect 5418 309922 5514 309978
rect 5570 309922 5638 309978
rect 5694 309922 5762 309978
rect 5818 309922 5886 309978
rect 5942 309922 6038 309978
rect -956 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 -336 292350
rect -956 292226 -336 292294
rect -956 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 -336 292226
rect -956 292102 -336 292170
rect -956 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 -336 292102
rect -956 291978 -336 292046
rect -956 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 -336 291978
rect -956 274350 -336 291922
rect 5418 292350 6038 309922
rect 12448 310350 12768 310384
rect 12448 310294 12518 310350
rect 12574 310294 12642 310350
rect 12698 310294 12768 310350
rect 12448 310226 12768 310294
rect 12448 310170 12518 310226
rect 12574 310170 12642 310226
rect 12698 310170 12768 310226
rect 12448 310102 12768 310170
rect 12448 310046 12518 310102
rect 12574 310046 12642 310102
rect 12698 310046 12768 310102
rect 12448 309978 12768 310046
rect 12448 309922 12518 309978
rect 12574 309922 12642 309978
rect 12698 309922 12768 309978
rect 12448 309888 12768 309922
rect 43168 310350 43488 310384
rect 43168 310294 43238 310350
rect 43294 310294 43362 310350
rect 43418 310294 43488 310350
rect 43168 310226 43488 310294
rect 43168 310170 43238 310226
rect 43294 310170 43362 310226
rect 43418 310170 43488 310226
rect 43168 310102 43488 310170
rect 43168 310046 43238 310102
rect 43294 310046 43362 310102
rect 43418 310046 43488 310102
rect 43168 309978 43488 310046
rect 43168 309922 43238 309978
rect 43294 309922 43362 309978
rect 43418 309922 43488 309978
rect 43168 309888 43488 309922
rect 73888 310350 74208 310384
rect 73888 310294 73958 310350
rect 74014 310294 74082 310350
rect 74138 310294 74208 310350
rect 73888 310226 74208 310294
rect 73888 310170 73958 310226
rect 74014 310170 74082 310226
rect 74138 310170 74208 310226
rect 73888 310102 74208 310170
rect 73888 310046 73958 310102
rect 74014 310046 74082 310102
rect 74138 310046 74208 310102
rect 73888 309978 74208 310046
rect 73888 309922 73958 309978
rect 74014 309922 74082 309978
rect 74138 309922 74208 309978
rect 73888 309888 74208 309922
rect 104608 310350 104928 310384
rect 104608 310294 104678 310350
rect 104734 310294 104802 310350
rect 104858 310294 104928 310350
rect 104608 310226 104928 310294
rect 104608 310170 104678 310226
rect 104734 310170 104802 310226
rect 104858 310170 104928 310226
rect 104608 310102 104928 310170
rect 104608 310046 104678 310102
rect 104734 310046 104802 310102
rect 104858 310046 104928 310102
rect 104608 309978 104928 310046
rect 104608 309922 104678 309978
rect 104734 309922 104802 309978
rect 104858 309922 104928 309978
rect 104608 309888 104928 309922
rect 135328 310350 135648 310384
rect 135328 310294 135398 310350
rect 135454 310294 135522 310350
rect 135578 310294 135648 310350
rect 135328 310226 135648 310294
rect 135328 310170 135398 310226
rect 135454 310170 135522 310226
rect 135578 310170 135648 310226
rect 135328 310102 135648 310170
rect 135328 310046 135398 310102
rect 135454 310046 135522 310102
rect 135578 310046 135648 310102
rect 135328 309978 135648 310046
rect 135328 309922 135398 309978
rect 135454 309922 135522 309978
rect 135578 309922 135648 309978
rect 135328 309888 135648 309922
rect 166048 310350 166368 310384
rect 166048 310294 166118 310350
rect 166174 310294 166242 310350
rect 166298 310294 166368 310350
rect 166048 310226 166368 310294
rect 166048 310170 166118 310226
rect 166174 310170 166242 310226
rect 166298 310170 166368 310226
rect 166048 310102 166368 310170
rect 166048 310046 166118 310102
rect 166174 310046 166242 310102
rect 166298 310046 166368 310102
rect 166048 309978 166368 310046
rect 166048 309922 166118 309978
rect 166174 309922 166242 309978
rect 166298 309922 166368 309978
rect 166048 309888 166368 309922
rect 196768 310350 197088 310384
rect 196768 310294 196838 310350
rect 196894 310294 196962 310350
rect 197018 310294 197088 310350
rect 196768 310226 197088 310294
rect 196768 310170 196838 310226
rect 196894 310170 196962 310226
rect 197018 310170 197088 310226
rect 196768 310102 197088 310170
rect 196768 310046 196838 310102
rect 196894 310046 196962 310102
rect 197018 310046 197088 310102
rect 196768 309978 197088 310046
rect 196768 309922 196838 309978
rect 196894 309922 196962 309978
rect 197018 309922 197088 309978
rect 196768 309888 197088 309922
rect 227488 310350 227808 310384
rect 227488 310294 227558 310350
rect 227614 310294 227682 310350
rect 227738 310294 227808 310350
rect 227488 310226 227808 310294
rect 227488 310170 227558 310226
rect 227614 310170 227682 310226
rect 227738 310170 227808 310226
rect 227488 310102 227808 310170
rect 227488 310046 227558 310102
rect 227614 310046 227682 310102
rect 227738 310046 227808 310102
rect 227488 309978 227808 310046
rect 227488 309922 227558 309978
rect 227614 309922 227682 309978
rect 227738 309922 227808 309978
rect 227488 309888 227808 309922
rect 258208 310350 258528 310384
rect 258208 310294 258278 310350
rect 258334 310294 258402 310350
rect 258458 310294 258528 310350
rect 258208 310226 258528 310294
rect 258208 310170 258278 310226
rect 258334 310170 258402 310226
rect 258458 310170 258528 310226
rect 258208 310102 258528 310170
rect 258208 310046 258278 310102
rect 258334 310046 258402 310102
rect 258458 310046 258528 310102
rect 258208 309978 258528 310046
rect 258208 309922 258278 309978
rect 258334 309922 258402 309978
rect 258458 309922 258528 309978
rect 258208 309888 258528 309922
rect 288928 310350 289248 310384
rect 288928 310294 288998 310350
rect 289054 310294 289122 310350
rect 289178 310294 289248 310350
rect 288928 310226 289248 310294
rect 288928 310170 288998 310226
rect 289054 310170 289122 310226
rect 289178 310170 289248 310226
rect 288928 310102 289248 310170
rect 288928 310046 288998 310102
rect 289054 310046 289122 310102
rect 289178 310046 289248 310102
rect 288928 309978 289248 310046
rect 288928 309922 288998 309978
rect 289054 309922 289122 309978
rect 289178 309922 289248 309978
rect 288928 309888 289248 309922
rect 319648 310350 319968 310384
rect 319648 310294 319718 310350
rect 319774 310294 319842 310350
rect 319898 310294 319968 310350
rect 319648 310226 319968 310294
rect 319648 310170 319718 310226
rect 319774 310170 319842 310226
rect 319898 310170 319968 310226
rect 319648 310102 319968 310170
rect 319648 310046 319718 310102
rect 319774 310046 319842 310102
rect 319898 310046 319968 310102
rect 319648 309978 319968 310046
rect 319648 309922 319718 309978
rect 319774 309922 319842 309978
rect 319898 309922 319968 309978
rect 319648 309888 319968 309922
rect 350368 310350 350688 310384
rect 350368 310294 350438 310350
rect 350494 310294 350562 310350
rect 350618 310294 350688 310350
rect 350368 310226 350688 310294
rect 350368 310170 350438 310226
rect 350494 310170 350562 310226
rect 350618 310170 350688 310226
rect 350368 310102 350688 310170
rect 350368 310046 350438 310102
rect 350494 310046 350562 310102
rect 350618 310046 350688 310102
rect 350368 309978 350688 310046
rect 350368 309922 350438 309978
rect 350494 309922 350562 309978
rect 350618 309922 350688 309978
rect 350368 309888 350688 309922
rect 381088 310350 381408 310384
rect 381088 310294 381158 310350
rect 381214 310294 381282 310350
rect 381338 310294 381408 310350
rect 381088 310226 381408 310294
rect 381088 310170 381158 310226
rect 381214 310170 381282 310226
rect 381338 310170 381408 310226
rect 381088 310102 381408 310170
rect 381088 310046 381158 310102
rect 381214 310046 381282 310102
rect 381338 310046 381408 310102
rect 381088 309978 381408 310046
rect 381088 309922 381158 309978
rect 381214 309922 381282 309978
rect 381338 309922 381408 309978
rect 381088 309888 381408 309922
rect 411808 310350 412128 310384
rect 411808 310294 411878 310350
rect 411934 310294 412002 310350
rect 412058 310294 412128 310350
rect 411808 310226 412128 310294
rect 411808 310170 411878 310226
rect 411934 310170 412002 310226
rect 412058 310170 412128 310226
rect 411808 310102 412128 310170
rect 411808 310046 411878 310102
rect 411934 310046 412002 310102
rect 412058 310046 412128 310102
rect 411808 309978 412128 310046
rect 411808 309922 411878 309978
rect 411934 309922 412002 309978
rect 412058 309922 412128 309978
rect 411808 309888 412128 309922
rect 442528 310350 442848 310384
rect 442528 310294 442598 310350
rect 442654 310294 442722 310350
rect 442778 310294 442848 310350
rect 442528 310226 442848 310294
rect 442528 310170 442598 310226
rect 442654 310170 442722 310226
rect 442778 310170 442848 310226
rect 442528 310102 442848 310170
rect 442528 310046 442598 310102
rect 442654 310046 442722 310102
rect 442778 310046 442848 310102
rect 442528 309978 442848 310046
rect 442528 309922 442598 309978
rect 442654 309922 442722 309978
rect 442778 309922 442848 309978
rect 442528 309888 442848 309922
rect 473248 310350 473568 310384
rect 473248 310294 473318 310350
rect 473374 310294 473442 310350
rect 473498 310294 473568 310350
rect 473248 310226 473568 310294
rect 473248 310170 473318 310226
rect 473374 310170 473442 310226
rect 473498 310170 473568 310226
rect 473248 310102 473568 310170
rect 473248 310046 473318 310102
rect 473374 310046 473442 310102
rect 473498 310046 473568 310102
rect 473248 309978 473568 310046
rect 473248 309922 473318 309978
rect 473374 309922 473442 309978
rect 473498 309922 473568 309978
rect 473248 309888 473568 309922
rect 503968 310350 504288 310384
rect 503968 310294 504038 310350
rect 504094 310294 504162 310350
rect 504218 310294 504288 310350
rect 503968 310226 504288 310294
rect 503968 310170 504038 310226
rect 504094 310170 504162 310226
rect 504218 310170 504288 310226
rect 503968 310102 504288 310170
rect 503968 310046 504038 310102
rect 504094 310046 504162 310102
rect 504218 310046 504288 310102
rect 503968 309978 504288 310046
rect 503968 309922 504038 309978
rect 504094 309922 504162 309978
rect 504218 309922 504288 309978
rect 503968 309888 504288 309922
rect 534688 310350 535008 310384
rect 534688 310294 534758 310350
rect 534814 310294 534882 310350
rect 534938 310294 535008 310350
rect 534688 310226 535008 310294
rect 534688 310170 534758 310226
rect 534814 310170 534882 310226
rect 534938 310170 535008 310226
rect 534688 310102 535008 310170
rect 534688 310046 534758 310102
rect 534814 310046 534882 310102
rect 534938 310046 535008 310102
rect 534688 309978 535008 310046
rect 534688 309922 534758 309978
rect 534814 309922 534882 309978
rect 534938 309922 535008 309978
rect 534688 309888 535008 309922
rect 565408 310350 565728 310384
rect 565408 310294 565478 310350
rect 565534 310294 565602 310350
rect 565658 310294 565728 310350
rect 565408 310226 565728 310294
rect 565408 310170 565478 310226
rect 565534 310170 565602 310226
rect 565658 310170 565728 310226
rect 565408 310102 565728 310170
rect 565408 310046 565478 310102
rect 565534 310046 565602 310102
rect 565658 310046 565728 310102
rect 565408 309978 565728 310046
rect 565408 309922 565478 309978
rect 565534 309922 565602 309978
rect 565658 309922 565728 309978
rect 565408 309888 565728 309922
rect 5418 292294 5514 292350
rect 5570 292294 5638 292350
rect 5694 292294 5762 292350
rect 5818 292294 5886 292350
rect 5942 292294 6038 292350
rect 5418 292226 6038 292294
rect 5418 292170 5514 292226
rect 5570 292170 5638 292226
rect 5694 292170 5762 292226
rect 5818 292170 5886 292226
rect 5942 292170 6038 292226
rect 5418 292102 6038 292170
rect 5418 292046 5514 292102
rect 5570 292046 5638 292102
rect 5694 292046 5762 292102
rect 5818 292046 5886 292102
rect 5942 292046 6038 292102
rect 5418 291978 6038 292046
rect 5418 291922 5514 291978
rect 5570 291922 5638 291978
rect 5694 291922 5762 291978
rect 5818 291922 5886 291978
rect 5942 291922 6038 291978
rect -956 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 -336 274350
rect -956 274226 -336 274294
rect -956 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 -336 274226
rect -956 274102 -336 274170
rect -956 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 -336 274102
rect -956 273978 -336 274046
rect -956 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 -336 273978
rect -956 256350 -336 273922
rect 4172 290836 4228 290846
rect 4172 270340 4228 290780
rect 4172 270274 4228 270284
rect 4284 276724 4340 276734
rect 4284 259812 4340 276668
rect 4284 259746 4340 259756
rect 5418 274350 6038 291922
rect 6188 304948 6244 304958
rect 6188 291396 6244 304892
rect 27808 298350 28128 298384
rect 27808 298294 27878 298350
rect 27934 298294 28002 298350
rect 28058 298294 28128 298350
rect 27808 298226 28128 298294
rect 27808 298170 27878 298226
rect 27934 298170 28002 298226
rect 28058 298170 28128 298226
rect 27808 298102 28128 298170
rect 27808 298046 27878 298102
rect 27934 298046 28002 298102
rect 28058 298046 28128 298102
rect 27808 297978 28128 298046
rect 27808 297922 27878 297978
rect 27934 297922 28002 297978
rect 28058 297922 28128 297978
rect 27808 297888 28128 297922
rect 58528 298350 58848 298384
rect 58528 298294 58598 298350
rect 58654 298294 58722 298350
rect 58778 298294 58848 298350
rect 58528 298226 58848 298294
rect 58528 298170 58598 298226
rect 58654 298170 58722 298226
rect 58778 298170 58848 298226
rect 58528 298102 58848 298170
rect 58528 298046 58598 298102
rect 58654 298046 58722 298102
rect 58778 298046 58848 298102
rect 58528 297978 58848 298046
rect 58528 297922 58598 297978
rect 58654 297922 58722 297978
rect 58778 297922 58848 297978
rect 58528 297888 58848 297922
rect 89248 298350 89568 298384
rect 89248 298294 89318 298350
rect 89374 298294 89442 298350
rect 89498 298294 89568 298350
rect 89248 298226 89568 298294
rect 89248 298170 89318 298226
rect 89374 298170 89442 298226
rect 89498 298170 89568 298226
rect 89248 298102 89568 298170
rect 89248 298046 89318 298102
rect 89374 298046 89442 298102
rect 89498 298046 89568 298102
rect 89248 297978 89568 298046
rect 89248 297922 89318 297978
rect 89374 297922 89442 297978
rect 89498 297922 89568 297978
rect 89248 297888 89568 297922
rect 119968 298350 120288 298384
rect 119968 298294 120038 298350
rect 120094 298294 120162 298350
rect 120218 298294 120288 298350
rect 119968 298226 120288 298294
rect 119968 298170 120038 298226
rect 120094 298170 120162 298226
rect 120218 298170 120288 298226
rect 119968 298102 120288 298170
rect 119968 298046 120038 298102
rect 120094 298046 120162 298102
rect 120218 298046 120288 298102
rect 119968 297978 120288 298046
rect 119968 297922 120038 297978
rect 120094 297922 120162 297978
rect 120218 297922 120288 297978
rect 119968 297888 120288 297922
rect 150688 298350 151008 298384
rect 150688 298294 150758 298350
rect 150814 298294 150882 298350
rect 150938 298294 151008 298350
rect 150688 298226 151008 298294
rect 150688 298170 150758 298226
rect 150814 298170 150882 298226
rect 150938 298170 151008 298226
rect 150688 298102 151008 298170
rect 150688 298046 150758 298102
rect 150814 298046 150882 298102
rect 150938 298046 151008 298102
rect 150688 297978 151008 298046
rect 150688 297922 150758 297978
rect 150814 297922 150882 297978
rect 150938 297922 151008 297978
rect 150688 297888 151008 297922
rect 181408 298350 181728 298384
rect 181408 298294 181478 298350
rect 181534 298294 181602 298350
rect 181658 298294 181728 298350
rect 181408 298226 181728 298294
rect 181408 298170 181478 298226
rect 181534 298170 181602 298226
rect 181658 298170 181728 298226
rect 181408 298102 181728 298170
rect 181408 298046 181478 298102
rect 181534 298046 181602 298102
rect 181658 298046 181728 298102
rect 181408 297978 181728 298046
rect 181408 297922 181478 297978
rect 181534 297922 181602 297978
rect 181658 297922 181728 297978
rect 181408 297888 181728 297922
rect 212128 298350 212448 298384
rect 212128 298294 212198 298350
rect 212254 298294 212322 298350
rect 212378 298294 212448 298350
rect 212128 298226 212448 298294
rect 212128 298170 212198 298226
rect 212254 298170 212322 298226
rect 212378 298170 212448 298226
rect 212128 298102 212448 298170
rect 212128 298046 212198 298102
rect 212254 298046 212322 298102
rect 212378 298046 212448 298102
rect 212128 297978 212448 298046
rect 212128 297922 212198 297978
rect 212254 297922 212322 297978
rect 212378 297922 212448 297978
rect 212128 297888 212448 297922
rect 242848 298350 243168 298384
rect 242848 298294 242918 298350
rect 242974 298294 243042 298350
rect 243098 298294 243168 298350
rect 242848 298226 243168 298294
rect 242848 298170 242918 298226
rect 242974 298170 243042 298226
rect 243098 298170 243168 298226
rect 242848 298102 243168 298170
rect 242848 298046 242918 298102
rect 242974 298046 243042 298102
rect 243098 298046 243168 298102
rect 242848 297978 243168 298046
rect 242848 297922 242918 297978
rect 242974 297922 243042 297978
rect 243098 297922 243168 297978
rect 242848 297888 243168 297922
rect 273568 298350 273888 298384
rect 273568 298294 273638 298350
rect 273694 298294 273762 298350
rect 273818 298294 273888 298350
rect 273568 298226 273888 298294
rect 273568 298170 273638 298226
rect 273694 298170 273762 298226
rect 273818 298170 273888 298226
rect 273568 298102 273888 298170
rect 273568 298046 273638 298102
rect 273694 298046 273762 298102
rect 273818 298046 273888 298102
rect 273568 297978 273888 298046
rect 273568 297922 273638 297978
rect 273694 297922 273762 297978
rect 273818 297922 273888 297978
rect 273568 297888 273888 297922
rect 304288 298350 304608 298384
rect 304288 298294 304358 298350
rect 304414 298294 304482 298350
rect 304538 298294 304608 298350
rect 304288 298226 304608 298294
rect 304288 298170 304358 298226
rect 304414 298170 304482 298226
rect 304538 298170 304608 298226
rect 304288 298102 304608 298170
rect 304288 298046 304358 298102
rect 304414 298046 304482 298102
rect 304538 298046 304608 298102
rect 304288 297978 304608 298046
rect 304288 297922 304358 297978
rect 304414 297922 304482 297978
rect 304538 297922 304608 297978
rect 304288 297888 304608 297922
rect 335008 298350 335328 298384
rect 335008 298294 335078 298350
rect 335134 298294 335202 298350
rect 335258 298294 335328 298350
rect 335008 298226 335328 298294
rect 335008 298170 335078 298226
rect 335134 298170 335202 298226
rect 335258 298170 335328 298226
rect 335008 298102 335328 298170
rect 335008 298046 335078 298102
rect 335134 298046 335202 298102
rect 335258 298046 335328 298102
rect 335008 297978 335328 298046
rect 335008 297922 335078 297978
rect 335134 297922 335202 297978
rect 335258 297922 335328 297978
rect 335008 297888 335328 297922
rect 365728 298350 366048 298384
rect 365728 298294 365798 298350
rect 365854 298294 365922 298350
rect 365978 298294 366048 298350
rect 365728 298226 366048 298294
rect 365728 298170 365798 298226
rect 365854 298170 365922 298226
rect 365978 298170 366048 298226
rect 365728 298102 366048 298170
rect 365728 298046 365798 298102
rect 365854 298046 365922 298102
rect 365978 298046 366048 298102
rect 365728 297978 366048 298046
rect 365728 297922 365798 297978
rect 365854 297922 365922 297978
rect 365978 297922 366048 297978
rect 365728 297888 366048 297922
rect 396448 298350 396768 298384
rect 396448 298294 396518 298350
rect 396574 298294 396642 298350
rect 396698 298294 396768 298350
rect 396448 298226 396768 298294
rect 396448 298170 396518 298226
rect 396574 298170 396642 298226
rect 396698 298170 396768 298226
rect 396448 298102 396768 298170
rect 396448 298046 396518 298102
rect 396574 298046 396642 298102
rect 396698 298046 396768 298102
rect 396448 297978 396768 298046
rect 396448 297922 396518 297978
rect 396574 297922 396642 297978
rect 396698 297922 396768 297978
rect 396448 297888 396768 297922
rect 427168 298350 427488 298384
rect 427168 298294 427238 298350
rect 427294 298294 427362 298350
rect 427418 298294 427488 298350
rect 427168 298226 427488 298294
rect 427168 298170 427238 298226
rect 427294 298170 427362 298226
rect 427418 298170 427488 298226
rect 427168 298102 427488 298170
rect 427168 298046 427238 298102
rect 427294 298046 427362 298102
rect 427418 298046 427488 298102
rect 427168 297978 427488 298046
rect 427168 297922 427238 297978
rect 427294 297922 427362 297978
rect 427418 297922 427488 297978
rect 427168 297888 427488 297922
rect 457888 298350 458208 298384
rect 457888 298294 457958 298350
rect 458014 298294 458082 298350
rect 458138 298294 458208 298350
rect 457888 298226 458208 298294
rect 457888 298170 457958 298226
rect 458014 298170 458082 298226
rect 458138 298170 458208 298226
rect 457888 298102 458208 298170
rect 457888 298046 457958 298102
rect 458014 298046 458082 298102
rect 458138 298046 458208 298102
rect 457888 297978 458208 298046
rect 457888 297922 457958 297978
rect 458014 297922 458082 297978
rect 458138 297922 458208 297978
rect 457888 297888 458208 297922
rect 488608 298350 488928 298384
rect 488608 298294 488678 298350
rect 488734 298294 488802 298350
rect 488858 298294 488928 298350
rect 488608 298226 488928 298294
rect 488608 298170 488678 298226
rect 488734 298170 488802 298226
rect 488858 298170 488928 298226
rect 488608 298102 488928 298170
rect 488608 298046 488678 298102
rect 488734 298046 488802 298102
rect 488858 298046 488928 298102
rect 488608 297978 488928 298046
rect 488608 297922 488678 297978
rect 488734 297922 488802 297978
rect 488858 297922 488928 297978
rect 488608 297888 488928 297922
rect 519328 298350 519648 298384
rect 519328 298294 519398 298350
rect 519454 298294 519522 298350
rect 519578 298294 519648 298350
rect 519328 298226 519648 298294
rect 519328 298170 519398 298226
rect 519454 298170 519522 298226
rect 519578 298170 519648 298226
rect 519328 298102 519648 298170
rect 519328 298046 519398 298102
rect 519454 298046 519522 298102
rect 519578 298046 519648 298102
rect 519328 297978 519648 298046
rect 519328 297922 519398 297978
rect 519454 297922 519522 297978
rect 519578 297922 519648 297978
rect 519328 297888 519648 297922
rect 550048 298350 550368 298384
rect 550048 298294 550118 298350
rect 550174 298294 550242 298350
rect 550298 298294 550368 298350
rect 550048 298226 550368 298294
rect 550048 298170 550118 298226
rect 550174 298170 550242 298226
rect 550298 298170 550368 298226
rect 550048 298102 550368 298170
rect 550048 298046 550118 298102
rect 550174 298046 550242 298102
rect 550298 298046 550368 298102
rect 550048 297978 550368 298046
rect 550048 297922 550118 297978
rect 550174 297922 550242 297978
rect 550298 297922 550368 297978
rect 550048 297888 550368 297922
rect 12448 292350 12768 292384
rect 12448 292294 12518 292350
rect 12574 292294 12642 292350
rect 12698 292294 12768 292350
rect 12448 292226 12768 292294
rect 12448 292170 12518 292226
rect 12574 292170 12642 292226
rect 12698 292170 12768 292226
rect 12448 292102 12768 292170
rect 12448 292046 12518 292102
rect 12574 292046 12642 292102
rect 12698 292046 12768 292102
rect 12448 291978 12768 292046
rect 12448 291922 12518 291978
rect 12574 291922 12642 291978
rect 12698 291922 12768 291978
rect 12448 291888 12768 291922
rect 43168 292350 43488 292384
rect 43168 292294 43238 292350
rect 43294 292294 43362 292350
rect 43418 292294 43488 292350
rect 43168 292226 43488 292294
rect 43168 292170 43238 292226
rect 43294 292170 43362 292226
rect 43418 292170 43488 292226
rect 43168 292102 43488 292170
rect 43168 292046 43238 292102
rect 43294 292046 43362 292102
rect 43418 292046 43488 292102
rect 43168 291978 43488 292046
rect 43168 291922 43238 291978
rect 43294 291922 43362 291978
rect 43418 291922 43488 291978
rect 43168 291888 43488 291922
rect 73888 292350 74208 292384
rect 73888 292294 73958 292350
rect 74014 292294 74082 292350
rect 74138 292294 74208 292350
rect 73888 292226 74208 292294
rect 73888 292170 73958 292226
rect 74014 292170 74082 292226
rect 74138 292170 74208 292226
rect 73888 292102 74208 292170
rect 73888 292046 73958 292102
rect 74014 292046 74082 292102
rect 74138 292046 74208 292102
rect 73888 291978 74208 292046
rect 73888 291922 73958 291978
rect 74014 291922 74082 291978
rect 74138 291922 74208 291978
rect 73888 291888 74208 291922
rect 104608 292350 104928 292384
rect 104608 292294 104678 292350
rect 104734 292294 104802 292350
rect 104858 292294 104928 292350
rect 104608 292226 104928 292294
rect 104608 292170 104678 292226
rect 104734 292170 104802 292226
rect 104858 292170 104928 292226
rect 104608 292102 104928 292170
rect 104608 292046 104678 292102
rect 104734 292046 104802 292102
rect 104858 292046 104928 292102
rect 104608 291978 104928 292046
rect 104608 291922 104678 291978
rect 104734 291922 104802 291978
rect 104858 291922 104928 291978
rect 104608 291888 104928 291922
rect 135328 292350 135648 292384
rect 135328 292294 135398 292350
rect 135454 292294 135522 292350
rect 135578 292294 135648 292350
rect 135328 292226 135648 292294
rect 135328 292170 135398 292226
rect 135454 292170 135522 292226
rect 135578 292170 135648 292226
rect 135328 292102 135648 292170
rect 135328 292046 135398 292102
rect 135454 292046 135522 292102
rect 135578 292046 135648 292102
rect 135328 291978 135648 292046
rect 135328 291922 135398 291978
rect 135454 291922 135522 291978
rect 135578 291922 135648 291978
rect 135328 291888 135648 291922
rect 166048 292350 166368 292384
rect 166048 292294 166118 292350
rect 166174 292294 166242 292350
rect 166298 292294 166368 292350
rect 166048 292226 166368 292294
rect 166048 292170 166118 292226
rect 166174 292170 166242 292226
rect 166298 292170 166368 292226
rect 166048 292102 166368 292170
rect 166048 292046 166118 292102
rect 166174 292046 166242 292102
rect 166298 292046 166368 292102
rect 166048 291978 166368 292046
rect 166048 291922 166118 291978
rect 166174 291922 166242 291978
rect 166298 291922 166368 291978
rect 166048 291888 166368 291922
rect 196768 292350 197088 292384
rect 196768 292294 196838 292350
rect 196894 292294 196962 292350
rect 197018 292294 197088 292350
rect 196768 292226 197088 292294
rect 196768 292170 196838 292226
rect 196894 292170 196962 292226
rect 197018 292170 197088 292226
rect 196768 292102 197088 292170
rect 196768 292046 196838 292102
rect 196894 292046 196962 292102
rect 197018 292046 197088 292102
rect 196768 291978 197088 292046
rect 196768 291922 196838 291978
rect 196894 291922 196962 291978
rect 197018 291922 197088 291978
rect 196768 291888 197088 291922
rect 227488 292350 227808 292384
rect 227488 292294 227558 292350
rect 227614 292294 227682 292350
rect 227738 292294 227808 292350
rect 227488 292226 227808 292294
rect 227488 292170 227558 292226
rect 227614 292170 227682 292226
rect 227738 292170 227808 292226
rect 227488 292102 227808 292170
rect 227488 292046 227558 292102
rect 227614 292046 227682 292102
rect 227738 292046 227808 292102
rect 227488 291978 227808 292046
rect 227488 291922 227558 291978
rect 227614 291922 227682 291978
rect 227738 291922 227808 291978
rect 227488 291888 227808 291922
rect 258208 292350 258528 292384
rect 258208 292294 258278 292350
rect 258334 292294 258402 292350
rect 258458 292294 258528 292350
rect 258208 292226 258528 292294
rect 258208 292170 258278 292226
rect 258334 292170 258402 292226
rect 258458 292170 258528 292226
rect 258208 292102 258528 292170
rect 258208 292046 258278 292102
rect 258334 292046 258402 292102
rect 258458 292046 258528 292102
rect 258208 291978 258528 292046
rect 258208 291922 258278 291978
rect 258334 291922 258402 291978
rect 258458 291922 258528 291978
rect 258208 291888 258528 291922
rect 288928 292350 289248 292384
rect 288928 292294 288998 292350
rect 289054 292294 289122 292350
rect 289178 292294 289248 292350
rect 288928 292226 289248 292294
rect 288928 292170 288998 292226
rect 289054 292170 289122 292226
rect 289178 292170 289248 292226
rect 288928 292102 289248 292170
rect 288928 292046 288998 292102
rect 289054 292046 289122 292102
rect 289178 292046 289248 292102
rect 288928 291978 289248 292046
rect 288928 291922 288998 291978
rect 289054 291922 289122 291978
rect 289178 291922 289248 291978
rect 288928 291888 289248 291922
rect 319648 292350 319968 292384
rect 319648 292294 319718 292350
rect 319774 292294 319842 292350
rect 319898 292294 319968 292350
rect 319648 292226 319968 292294
rect 319648 292170 319718 292226
rect 319774 292170 319842 292226
rect 319898 292170 319968 292226
rect 319648 292102 319968 292170
rect 319648 292046 319718 292102
rect 319774 292046 319842 292102
rect 319898 292046 319968 292102
rect 319648 291978 319968 292046
rect 319648 291922 319718 291978
rect 319774 291922 319842 291978
rect 319898 291922 319968 291978
rect 319648 291888 319968 291922
rect 350368 292350 350688 292384
rect 350368 292294 350438 292350
rect 350494 292294 350562 292350
rect 350618 292294 350688 292350
rect 350368 292226 350688 292294
rect 350368 292170 350438 292226
rect 350494 292170 350562 292226
rect 350618 292170 350688 292226
rect 350368 292102 350688 292170
rect 350368 292046 350438 292102
rect 350494 292046 350562 292102
rect 350618 292046 350688 292102
rect 350368 291978 350688 292046
rect 350368 291922 350438 291978
rect 350494 291922 350562 291978
rect 350618 291922 350688 291978
rect 350368 291888 350688 291922
rect 381088 292350 381408 292384
rect 381088 292294 381158 292350
rect 381214 292294 381282 292350
rect 381338 292294 381408 292350
rect 381088 292226 381408 292294
rect 381088 292170 381158 292226
rect 381214 292170 381282 292226
rect 381338 292170 381408 292226
rect 381088 292102 381408 292170
rect 381088 292046 381158 292102
rect 381214 292046 381282 292102
rect 381338 292046 381408 292102
rect 381088 291978 381408 292046
rect 381088 291922 381158 291978
rect 381214 291922 381282 291978
rect 381338 291922 381408 291978
rect 381088 291888 381408 291922
rect 411808 292350 412128 292384
rect 411808 292294 411878 292350
rect 411934 292294 412002 292350
rect 412058 292294 412128 292350
rect 411808 292226 412128 292294
rect 411808 292170 411878 292226
rect 411934 292170 412002 292226
rect 412058 292170 412128 292226
rect 411808 292102 412128 292170
rect 411808 292046 411878 292102
rect 411934 292046 412002 292102
rect 412058 292046 412128 292102
rect 411808 291978 412128 292046
rect 411808 291922 411878 291978
rect 411934 291922 412002 291978
rect 412058 291922 412128 291978
rect 411808 291888 412128 291922
rect 442528 292350 442848 292384
rect 442528 292294 442598 292350
rect 442654 292294 442722 292350
rect 442778 292294 442848 292350
rect 442528 292226 442848 292294
rect 442528 292170 442598 292226
rect 442654 292170 442722 292226
rect 442778 292170 442848 292226
rect 442528 292102 442848 292170
rect 442528 292046 442598 292102
rect 442654 292046 442722 292102
rect 442778 292046 442848 292102
rect 442528 291978 442848 292046
rect 442528 291922 442598 291978
rect 442654 291922 442722 291978
rect 442778 291922 442848 291978
rect 442528 291888 442848 291922
rect 473248 292350 473568 292384
rect 473248 292294 473318 292350
rect 473374 292294 473442 292350
rect 473498 292294 473568 292350
rect 473248 292226 473568 292294
rect 473248 292170 473318 292226
rect 473374 292170 473442 292226
rect 473498 292170 473568 292226
rect 473248 292102 473568 292170
rect 473248 292046 473318 292102
rect 473374 292046 473442 292102
rect 473498 292046 473568 292102
rect 473248 291978 473568 292046
rect 473248 291922 473318 291978
rect 473374 291922 473442 291978
rect 473498 291922 473568 291978
rect 473248 291888 473568 291922
rect 503968 292350 504288 292384
rect 503968 292294 504038 292350
rect 504094 292294 504162 292350
rect 504218 292294 504288 292350
rect 503968 292226 504288 292294
rect 503968 292170 504038 292226
rect 504094 292170 504162 292226
rect 504218 292170 504288 292226
rect 503968 292102 504288 292170
rect 503968 292046 504038 292102
rect 504094 292046 504162 292102
rect 504218 292046 504288 292102
rect 503968 291978 504288 292046
rect 503968 291922 504038 291978
rect 504094 291922 504162 291978
rect 504218 291922 504288 291978
rect 503968 291888 504288 291922
rect 534688 292350 535008 292384
rect 534688 292294 534758 292350
rect 534814 292294 534882 292350
rect 534938 292294 535008 292350
rect 534688 292226 535008 292294
rect 534688 292170 534758 292226
rect 534814 292170 534882 292226
rect 534938 292170 535008 292226
rect 534688 292102 535008 292170
rect 534688 292046 534758 292102
rect 534814 292046 534882 292102
rect 534938 292046 535008 292102
rect 534688 291978 535008 292046
rect 534688 291922 534758 291978
rect 534814 291922 534882 291978
rect 534938 291922 535008 291978
rect 534688 291888 535008 291922
rect 565408 292350 565728 292384
rect 565408 292294 565478 292350
rect 565534 292294 565602 292350
rect 565658 292294 565728 292350
rect 565408 292226 565728 292294
rect 565408 292170 565478 292226
rect 565534 292170 565602 292226
rect 565658 292170 565728 292226
rect 565408 292102 565728 292170
rect 565408 292046 565478 292102
rect 565534 292046 565602 292102
rect 565658 292046 565728 292102
rect 565408 291978 565728 292046
rect 565408 291922 565478 291978
rect 565534 291922 565602 291978
rect 565658 291922 565728 291978
rect 565408 291888 565728 291922
rect 6188 291330 6244 291340
rect 27808 280350 28128 280384
rect 27808 280294 27878 280350
rect 27934 280294 28002 280350
rect 28058 280294 28128 280350
rect 27808 280226 28128 280294
rect 27808 280170 27878 280226
rect 27934 280170 28002 280226
rect 28058 280170 28128 280226
rect 27808 280102 28128 280170
rect 27808 280046 27878 280102
rect 27934 280046 28002 280102
rect 28058 280046 28128 280102
rect 27808 279978 28128 280046
rect 27808 279922 27878 279978
rect 27934 279922 28002 279978
rect 28058 279922 28128 279978
rect 27808 279888 28128 279922
rect 58528 280350 58848 280384
rect 58528 280294 58598 280350
rect 58654 280294 58722 280350
rect 58778 280294 58848 280350
rect 58528 280226 58848 280294
rect 58528 280170 58598 280226
rect 58654 280170 58722 280226
rect 58778 280170 58848 280226
rect 58528 280102 58848 280170
rect 58528 280046 58598 280102
rect 58654 280046 58722 280102
rect 58778 280046 58848 280102
rect 58528 279978 58848 280046
rect 58528 279922 58598 279978
rect 58654 279922 58722 279978
rect 58778 279922 58848 279978
rect 58528 279888 58848 279922
rect 89248 280350 89568 280384
rect 89248 280294 89318 280350
rect 89374 280294 89442 280350
rect 89498 280294 89568 280350
rect 89248 280226 89568 280294
rect 89248 280170 89318 280226
rect 89374 280170 89442 280226
rect 89498 280170 89568 280226
rect 89248 280102 89568 280170
rect 89248 280046 89318 280102
rect 89374 280046 89442 280102
rect 89498 280046 89568 280102
rect 89248 279978 89568 280046
rect 89248 279922 89318 279978
rect 89374 279922 89442 279978
rect 89498 279922 89568 279978
rect 89248 279888 89568 279922
rect 119968 280350 120288 280384
rect 119968 280294 120038 280350
rect 120094 280294 120162 280350
rect 120218 280294 120288 280350
rect 119968 280226 120288 280294
rect 119968 280170 120038 280226
rect 120094 280170 120162 280226
rect 120218 280170 120288 280226
rect 119968 280102 120288 280170
rect 119968 280046 120038 280102
rect 120094 280046 120162 280102
rect 120218 280046 120288 280102
rect 119968 279978 120288 280046
rect 119968 279922 120038 279978
rect 120094 279922 120162 279978
rect 120218 279922 120288 279978
rect 119968 279888 120288 279922
rect 150688 280350 151008 280384
rect 150688 280294 150758 280350
rect 150814 280294 150882 280350
rect 150938 280294 151008 280350
rect 150688 280226 151008 280294
rect 150688 280170 150758 280226
rect 150814 280170 150882 280226
rect 150938 280170 151008 280226
rect 150688 280102 151008 280170
rect 150688 280046 150758 280102
rect 150814 280046 150882 280102
rect 150938 280046 151008 280102
rect 150688 279978 151008 280046
rect 150688 279922 150758 279978
rect 150814 279922 150882 279978
rect 150938 279922 151008 279978
rect 150688 279888 151008 279922
rect 181408 280350 181728 280384
rect 181408 280294 181478 280350
rect 181534 280294 181602 280350
rect 181658 280294 181728 280350
rect 181408 280226 181728 280294
rect 181408 280170 181478 280226
rect 181534 280170 181602 280226
rect 181658 280170 181728 280226
rect 181408 280102 181728 280170
rect 181408 280046 181478 280102
rect 181534 280046 181602 280102
rect 181658 280046 181728 280102
rect 181408 279978 181728 280046
rect 181408 279922 181478 279978
rect 181534 279922 181602 279978
rect 181658 279922 181728 279978
rect 181408 279888 181728 279922
rect 212128 280350 212448 280384
rect 212128 280294 212198 280350
rect 212254 280294 212322 280350
rect 212378 280294 212448 280350
rect 212128 280226 212448 280294
rect 212128 280170 212198 280226
rect 212254 280170 212322 280226
rect 212378 280170 212448 280226
rect 212128 280102 212448 280170
rect 212128 280046 212198 280102
rect 212254 280046 212322 280102
rect 212378 280046 212448 280102
rect 212128 279978 212448 280046
rect 212128 279922 212198 279978
rect 212254 279922 212322 279978
rect 212378 279922 212448 279978
rect 212128 279888 212448 279922
rect 242848 280350 243168 280384
rect 242848 280294 242918 280350
rect 242974 280294 243042 280350
rect 243098 280294 243168 280350
rect 242848 280226 243168 280294
rect 242848 280170 242918 280226
rect 242974 280170 243042 280226
rect 243098 280170 243168 280226
rect 242848 280102 243168 280170
rect 242848 280046 242918 280102
rect 242974 280046 243042 280102
rect 243098 280046 243168 280102
rect 242848 279978 243168 280046
rect 242848 279922 242918 279978
rect 242974 279922 243042 279978
rect 243098 279922 243168 279978
rect 242848 279888 243168 279922
rect 273568 280350 273888 280384
rect 273568 280294 273638 280350
rect 273694 280294 273762 280350
rect 273818 280294 273888 280350
rect 273568 280226 273888 280294
rect 273568 280170 273638 280226
rect 273694 280170 273762 280226
rect 273818 280170 273888 280226
rect 273568 280102 273888 280170
rect 273568 280046 273638 280102
rect 273694 280046 273762 280102
rect 273818 280046 273888 280102
rect 273568 279978 273888 280046
rect 273568 279922 273638 279978
rect 273694 279922 273762 279978
rect 273818 279922 273888 279978
rect 273568 279888 273888 279922
rect 304288 280350 304608 280384
rect 304288 280294 304358 280350
rect 304414 280294 304482 280350
rect 304538 280294 304608 280350
rect 304288 280226 304608 280294
rect 304288 280170 304358 280226
rect 304414 280170 304482 280226
rect 304538 280170 304608 280226
rect 304288 280102 304608 280170
rect 304288 280046 304358 280102
rect 304414 280046 304482 280102
rect 304538 280046 304608 280102
rect 304288 279978 304608 280046
rect 304288 279922 304358 279978
rect 304414 279922 304482 279978
rect 304538 279922 304608 279978
rect 304288 279888 304608 279922
rect 335008 280350 335328 280384
rect 335008 280294 335078 280350
rect 335134 280294 335202 280350
rect 335258 280294 335328 280350
rect 335008 280226 335328 280294
rect 335008 280170 335078 280226
rect 335134 280170 335202 280226
rect 335258 280170 335328 280226
rect 335008 280102 335328 280170
rect 335008 280046 335078 280102
rect 335134 280046 335202 280102
rect 335258 280046 335328 280102
rect 335008 279978 335328 280046
rect 335008 279922 335078 279978
rect 335134 279922 335202 279978
rect 335258 279922 335328 279978
rect 335008 279888 335328 279922
rect 365728 280350 366048 280384
rect 365728 280294 365798 280350
rect 365854 280294 365922 280350
rect 365978 280294 366048 280350
rect 365728 280226 366048 280294
rect 365728 280170 365798 280226
rect 365854 280170 365922 280226
rect 365978 280170 366048 280226
rect 365728 280102 366048 280170
rect 365728 280046 365798 280102
rect 365854 280046 365922 280102
rect 365978 280046 366048 280102
rect 365728 279978 366048 280046
rect 365728 279922 365798 279978
rect 365854 279922 365922 279978
rect 365978 279922 366048 279978
rect 365728 279888 366048 279922
rect 396448 280350 396768 280384
rect 396448 280294 396518 280350
rect 396574 280294 396642 280350
rect 396698 280294 396768 280350
rect 396448 280226 396768 280294
rect 396448 280170 396518 280226
rect 396574 280170 396642 280226
rect 396698 280170 396768 280226
rect 396448 280102 396768 280170
rect 396448 280046 396518 280102
rect 396574 280046 396642 280102
rect 396698 280046 396768 280102
rect 396448 279978 396768 280046
rect 396448 279922 396518 279978
rect 396574 279922 396642 279978
rect 396698 279922 396768 279978
rect 396448 279888 396768 279922
rect 427168 280350 427488 280384
rect 427168 280294 427238 280350
rect 427294 280294 427362 280350
rect 427418 280294 427488 280350
rect 427168 280226 427488 280294
rect 427168 280170 427238 280226
rect 427294 280170 427362 280226
rect 427418 280170 427488 280226
rect 427168 280102 427488 280170
rect 427168 280046 427238 280102
rect 427294 280046 427362 280102
rect 427418 280046 427488 280102
rect 427168 279978 427488 280046
rect 427168 279922 427238 279978
rect 427294 279922 427362 279978
rect 427418 279922 427488 279978
rect 427168 279888 427488 279922
rect 457888 280350 458208 280384
rect 457888 280294 457958 280350
rect 458014 280294 458082 280350
rect 458138 280294 458208 280350
rect 457888 280226 458208 280294
rect 457888 280170 457958 280226
rect 458014 280170 458082 280226
rect 458138 280170 458208 280226
rect 457888 280102 458208 280170
rect 457888 280046 457958 280102
rect 458014 280046 458082 280102
rect 458138 280046 458208 280102
rect 457888 279978 458208 280046
rect 457888 279922 457958 279978
rect 458014 279922 458082 279978
rect 458138 279922 458208 279978
rect 457888 279888 458208 279922
rect 488608 280350 488928 280384
rect 488608 280294 488678 280350
rect 488734 280294 488802 280350
rect 488858 280294 488928 280350
rect 488608 280226 488928 280294
rect 488608 280170 488678 280226
rect 488734 280170 488802 280226
rect 488858 280170 488928 280226
rect 488608 280102 488928 280170
rect 488608 280046 488678 280102
rect 488734 280046 488802 280102
rect 488858 280046 488928 280102
rect 488608 279978 488928 280046
rect 488608 279922 488678 279978
rect 488734 279922 488802 279978
rect 488858 279922 488928 279978
rect 488608 279888 488928 279922
rect 519328 280350 519648 280384
rect 519328 280294 519398 280350
rect 519454 280294 519522 280350
rect 519578 280294 519648 280350
rect 519328 280226 519648 280294
rect 519328 280170 519398 280226
rect 519454 280170 519522 280226
rect 519578 280170 519648 280226
rect 519328 280102 519648 280170
rect 519328 280046 519398 280102
rect 519454 280046 519522 280102
rect 519578 280046 519648 280102
rect 519328 279978 519648 280046
rect 519328 279922 519398 279978
rect 519454 279922 519522 279978
rect 519578 279922 519648 279978
rect 519328 279888 519648 279922
rect 550048 280350 550368 280384
rect 550048 280294 550118 280350
rect 550174 280294 550242 280350
rect 550298 280294 550368 280350
rect 550048 280226 550368 280294
rect 550048 280170 550118 280226
rect 550174 280170 550242 280226
rect 550298 280170 550368 280226
rect 550048 280102 550368 280170
rect 550048 280046 550118 280102
rect 550174 280046 550242 280102
rect 550298 280046 550368 280102
rect 550048 279978 550368 280046
rect 550048 279922 550118 279978
rect 550174 279922 550242 279978
rect 550298 279922 550368 279978
rect 550048 279888 550368 279922
rect 585452 275268 585508 311052
rect 585564 296772 585620 324268
rect 585676 307524 585732 337484
rect 585676 307458 585732 307468
rect 589098 328350 589718 345922
rect 590492 363972 590548 363982
rect 590492 339780 590548 363916
rect 590492 339714 590548 339724
rect 592818 352350 593438 369922
rect 592818 352294 592914 352350
rect 592970 352294 593038 352350
rect 593094 352294 593162 352350
rect 593218 352294 593286 352350
rect 593342 352294 593438 352350
rect 592818 352226 593438 352294
rect 592818 352170 592914 352226
rect 592970 352170 593038 352226
rect 593094 352170 593162 352226
rect 593218 352170 593286 352226
rect 593342 352170 593438 352226
rect 592818 352102 593438 352170
rect 592818 352046 592914 352102
rect 592970 352046 593038 352102
rect 593094 352046 593162 352102
rect 593218 352046 593286 352102
rect 593342 352046 593438 352102
rect 592818 351978 593438 352046
rect 592818 351922 592914 351978
rect 592970 351922 593038 351978
rect 593094 351922 593162 351978
rect 593218 351922 593286 351978
rect 593342 351922 593438 351978
rect 589098 328294 589194 328350
rect 589250 328294 589318 328350
rect 589374 328294 589442 328350
rect 589498 328294 589566 328350
rect 589622 328294 589718 328350
rect 589098 328226 589718 328294
rect 589098 328170 589194 328226
rect 589250 328170 589318 328226
rect 589374 328170 589442 328226
rect 589498 328170 589566 328226
rect 589622 328170 589718 328226
rect 589098 328102 589718 328170
rect 589098 328046 589194 328102
rect 589250 328046 589318 328102
rect 589374 328046 589442 328102
rect 589498 328046 589566 328102
rect 589622 328046 589718 328102
rect 589098 327978 589718 328046
rect 589098 327922 589194 327978
rect 589250 327922 589318 327978
rect 589374 327922 589442 327978
rect 589498 327922 589566 327978
rect 589622 327922 589718 327978
rect 589098 310350 589718 327922
rect 589098 310294 589194 310350
rect 589250 310294 589318 310350
rect 589374 310294 589442 310350
rect 589498 310294 589566 310350
rect 589622 310294 589718 310350
rect 589098 310226 589718 310294
rect 589098 310170 589194 310226
rect 589250 310170 589318 310226
rect 589374 310170 589442 310226
rect 589498 310170 589566 310226
rect 589622 310170 589718 310226
rect 589098 310102 589718 310170
rect 589098 310046 589194 310102
rect 589250 310046 589318 310102
rect 589374 310046 589442 310102
rect 589498 310046 589566 310102
rect 589622 310046 589718 310102
rect 589098 309978 589718 310046
rect 589098 309922 589194 309978
rect 589250 309922 589318 309978
rect 589374 309922 589442 309978
rect 589498 309922 589566 309978
rect 589622 309922 589718 309978
rect 585564 296706 585620 296716
rect 589098 292350 589718 309922
rect 592818 334350 593438 351922
rect 592818 334294 592914 334350
rect 592970 334294 593038 334350
rect 593094 334294 593162 334350
rect 593218 334294 593286 334350
rect 593342 334294 593438 334350
rect 592818 334226 593438 334294
rect 592818 334170 592914 334226
rect 592970 334170 593038 334226
rect 593094 334170 593162 334226
rect 593218 334170 593286 334226
rect 593342 334170 593438 334226
rect 592818 334102 593438 334170
rect 592818 334046 592914 334102
rect 592970 334046 593038 334102
rect 593094 334046 593162 334102
rect 593218 334046 593286 334102
rect 593342 334046 593438 334102
rect 592818 333978 593438 334046
rect 592818 333922 592914 333978
rect 592970 333922 593038 333978
rect 593094 333922 593162 333978
rect 593218 333922 593286 333978
rect 593342 333922 593438 333978
rect 592818 316350 593438 333922
rect 592818 316294 592914 316350
rect 592970 316294 593038 316350
rect 593094 316294 593162 316350
rect 593218 316294 593286 316350
rect 593342 316294 593438 316350
rect 592818 316226 593438 316294
rect 592818 316170 592914 316226
rect 592970 316170 593038 316226
rect 593094 316170 593162 316226
rect 593218 316170 593286 316226
rect 593342 316170 593438 316226
rect 592818 316102 593438 316170
rect 592818 316046 592914 316102
rect 592970 316046 593038 316102
rect 593094 316046 593162 316102
rect 593218 316046 593286 316102
rect 593342 316046 593438 316102
rect 592818 315978 593438 316046
rect 592818 315922 592914 315978
rect 592970 315922 593038 315978
rect 593094 315922 593162 315978
rect 593218 315922 593286 315978
rect 593342 315922 593438 315978
rect 592818 298350 593438 315922
rect 592818 298294 592914 298350
rect 592970 298294 593038 298350
rect 593094 298294 593162 298350
rect 593218 298294 593286 298350
rect 593342 298294 593438 298350
rect 592818 298226 593438 298294
rect 592818 298170 592914 298226
rect 592970 298170 593038 298226
rect 593094 298170 593162 298226
rect 593218 298170 593286 298226
rect 593342 298170 593438 298226
rect 592818 298102 593438 298170
rect 592818 298046 592914 298102
rect 592970 298046 593038 298102
rect 593094 298046 593162 298102
rect 593218 298046 593286 298102
rect 593342 298046 593438 298102
rect 592818 297978 593438 298046
rect 592818 297922 592914 297978
rect 592970 297922 593038 297978
rect 593094 297922 593162 297978
rect 593218 297922 593286 297978
rect 593342 297922 593438 297978
rect 589098 292294 589194 292350
rect 589250 292294 589318 292350
rect 589374 292294 589442 292350
rect 589498 292294 589566 292350
rect 589622 292294 589718 292350
rect 589098 292226 589718 292294
rect 589098 292170 589194 292226
rect 589250 292170 589318 292226
rect 589374 292170 589442 292226
rect 589498 292170 589566 292226
rect 589622 292170 589718 292226
rect 589098 292102 589718 292170
rect 589098 292046 589194 292102
rect 589250 292046 589318 292102
rect 589374 292046 589442 292102
rect 589498 292046 589566 292102
rect 589622 292046 589718 292102
rect 589098 291978 589718 292046
rect 589098 291922 589194 291978
rect 589250 291922 589318 291978
rect 589374 291922 589442 291978
rect 589498 291922 589566 291978
rect 589622 291922 589718 291978
rect 585452 275202 585508 275212
rect 585564 284676 585620 284686
rect 5418 274294 5514 274350
rect 5570 274294 5638 274350
rect 5694 274294 5762 274350
rect 5818 274294 5886 274350
rect 5942 274294 6038 274350
rect 5418 274226 6038 274294
rect 5418 274170 5514 274226
rect 5570 274170 5638 274226
rect 5694 274170 5762 274226
rect 5818 274170 5886 274226
rect 5942 274170 6038 274226
rect 5418 274102 6038 274170
rect 5418 274046 5514 274102
rect 5570 274046 5638 274102
rect 5694 274046 5762 274102
rect 5818 274046 5886 274102
rect 5942 274046 6038 274102
rect 5418 273978 6038 274046
rect 5418 273922 5514 273978
rect 5570 273922 5638 273978
rect 5694 273922 5762 273978
rect 5818 273922 5886 273978
rect 5942 273922 6038 273978
rect -956 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 -336 256350
rect -956 256226 -336 256294
rect -956 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 -336 256226
rect -956 256102 -336 256170
rect -956 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 -336 256102
rect -956 255978 -336 256046
rect -956 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 -336 255978
rect -956 238350 -336 255922
rect -956 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 -336 238350
rect -956 238226 -336 238294
rect -956 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 -336 238226
rect -956 238102 -336 238170
rect -956 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 -336 238102
rect -956 237978 -336 238046
rect -956 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 -336 237978
rect -956 220350 -336 237922
rect 5418 256350 6038 273922
rect 12448 274350 12768 274384
rect 12448 274294 12518 274350
rect 12574 274294 12642 274350
rect 12698 274294 12768 274350
rect 12448 274226 12768 274294
rect 12448 274170 12518 274226
rect 12574 274170 12642 274226
rect 12698 274170 12768 274226
rect 12448 274102 12768 274170
rect 12448 274046 12518 274102
rect 12574 274046 12642 274102
rect 12698 274046 12768 274102
rect 12448 273978 12768 274046
rect 12448 273922 12518 273978
rect 12574 273922 12642 273978
rect 12698 273922 12768 273978
rect 12448 273888 12768 273922
rect 43168 274350 43488 274384
rect 43168 274294 43238 274350
rect 43294 274294 43362 274350
rect 43418 274294 43488 274350
rect 43168 274226 43488 274294
rect 43168 274170 43238 274226
rect 43294 274170 43362 274226
rect 43418 274170 43488 274226
rect 43168 274102 43488 274170
rect 43168 274046 43238 274102
rect 43294 274046 43362 274102
rect 43418 274046 43488 274102
rect 43168 273978 43488 274046
rect 43168 273922 43238 273978
rect 43294 273922 43362 273978
rect 43418 273922 43488 273978
rect 43168 273888 43488 273922
rect 73888 274350 74208 274384
rect 73888 274294 73958 274350
rect 74014 274294 74082 274350
rect 74138 274294 74208 274350
rect 73888 274226 74208 274294
rect 73888 274170 73958 274226
rect 74014 274170 74082 274226
rect 74138 274170 74208 274226
rect 73888 274102 74208 274170
rect 73888 274046 73958 274102
rect 74014 274046 74082 274102
rect 74138 274046 74208 274102
rect 73888 273978 74208 274046
rect 73888 273922 73958 273978
rect 74014 273922 74082 273978
rect 74138 273922 74208 273978
rect 73888 273888 74208 273922
rect 104608 274350 104928 274384
rect 104608 274294 104678 274350
rect 104734 274294 104802 274350
rect 104858 274294 104928 274350
rect 104608 274226 104928 274294
rect 104608 274170 104678 274226
rect 104734 274170 104802 274226
rect 104858 274170 104928 274226
rect 104608 274102 104928 274170
rect 104608 274046 104678 274102
rect 104734 274046 104802 274102
rect 104858 274046 104928 274102
rect 104608 273978 104928 274046
rect 104608 273922 104678 273978
rect 104734 273922 104802 273978
rect 104858 273922 104928 273978
rect 104608 273888 104928 273922
rect 135328 274350 135648 274384
rect 135328 274294 135398 274350
rect 135454 274294 135522 274350
rect 135578 274294 135648 274350
rect 135328 274226 135648 274294
rect 135328 274170 135398 274226
rect 135454 274170 135522 274226
rect 135578 274170 135648 274226
rect 135328 274102 135648 274170
rect 135328 274046 135398 274102
rect 135454 274046 135522 274102
rect 135578 274046 135648 274102
rect 135328 273978 135648 274046
rect 135328 273922 135398 273978
rect 135454 273922 135522 273978
rect 135578 273922 135648 273978
rect 135328 273888 135648 273922
rect 166048 274350 166368 274384
rect 166048 274294 166118 274350
rect 166174 274294 166242 274350
rect 166298 274294 166368 274350
rect 166048 274226 166368 274294
rect 166048 274170 166118 274226
rect 166174 274170 166242 274226
rect 166298 274170 166368 274226
rect 166048 274102 166368 274170
rect 166048 274046 166118 274102
rect 166174 274046 166242 274102
rect 166298 274046 166368 274102
rect 166048 273978 166368 274046
rect 166048 273922 166118 273978
rect 166174 273922 166242 273978
rect 166298 273922 166368 273978
rect 166048 273888 166368 273922
rect 196768 274350 197088 274384
rect 196768 274294 196838 274350
rect 196894 274294 196962 274350
rect 197018 274294 197088 274350
rect 196768 274226 197088 274294
rect 196768 274170 196838 274226
rect 196894 274170 196962 274226
rect 197018 274170 197088 274226
rect 196768 274102 197088 274170
rect 196768 274046 196838 274102
rect 196894 274046 196962 274102
rect 197018 274046 197088 274102
rect 196768 273978 197088 274046
rect 196768 273922 196838 273978
rect 196894 273922 196962 273978
rect 197018 273922 197088 273978
rect 196768 273888 197088 273922
rect 227488 274350 227808 274384
rect 227488 274294 227558 274350
rect 227614 274294 227682 274350
rect 227738 274294 227808 274350
rect 227488 274226 227808 274294
rect 227488 274170 227558 274226
rect 227614 274170 227682 274226
rect 227738 274170 227808 274226
rect 227488 274102 227808 274170
rect 227488 274046 227558 274102
rect 227614 274046 227682 274102
rect 227738 274046 227808 274102
rect 227488 273978 227808 274046
rect 227488 273922 227558 273978
rect 227614 273922 227682 273978
rect 227738 273922 227808 273978
rect 227488 273888 227808 273922
rect 258208 274350 258528 274384
rect 258208 274294 258278 274350
rect 258334 274294 258402 274350
rect 258458 274294 258528 274350
rect 258208 274226 258528 274294
rect 258208 274170 258278 274226
rect 258334 274170 258402 274226
rect 258458 274170 258528 274226
rect 258208 274102 258528 274170
rect 258208 274046 258278 274102
rect 258334 274046 258402 274102
rect 258458 274046 258528 274102
rect 258208 273978 258528 274046
rect 258208 273922 258278 273978
rect 258334 273922 258402 273978
rect 258458 273922 258528 273978
rect 258208 273888 258528 273922
rect 288928 274350 289248 274384
rect 288928 274294 288998 274350
rect 289054 274294 289122 274350
rect 289178 274294 289248 274350
rect 288928 274226 289248 274294
rect 288928 274170 288998 274226
rect 289054 274170 289122 274226
rect 289178 274170 289248 274226
rect 288928 274102 289248 274170
rect 288928 274046 288998 274102
rect 289054 274046 289122 274102
rect 289178 274046 289248 274102
rect 288928 273978 289248 274046
rect 288928 273922 288998 273978
rect 289054 273922 289122 273978
rect 289178 273922 289248 273978
rect 288928 273888 289248 273922
rect 319648 274350 319968 274384
rect 319648 274294 319718 274350
rect 319774 274294 319842 274350
rect 319898 274294 319968 274350
rect 319648 274226 319968 274294
rect 319648 274170 319718 274226
rect 319774 274170 319842 274226
rect 319898 274170 319968 274226
rect 319648 274102 319968 274170
rect 319648 274046 319718 274102
rect 319774 274046 319842 274102
rect 319898 274046 319968 274102
rect 319648 273978 319968 274046
rect 319648 273922 319718 273978
rect 319774 273922 319842 273978
rect 319898 273922 319968 273978
rect 319648 273888 319968 273922
rect 350368 274350 350688 274384
rect 350368 274294 350438 274350
rect 350494 274294 350562 274350
rect 350618 274294 350688 274350
rect 350368 274226 350688 274294
rect 350368 274170 350438 274226
rect 350494 274170 350562 274226
rect 350618 274170 350688 274226
rect 350368 274102 350688 274170
rect 350368 274046 350438 274102
rect 350494 274046 350562 274102
rect 350618 274046 350688 274102
rect 350368 273978 350688 274046
rect 350368 273922 350438 273978
rect 350494 273922 350562 273978
rect 350618 273922 350688 273978
rect 350368 273888 350688 273922
rect 381088 274350 381408 274384
rect 381088 274294 381158 274350
rect 381214 274294 381282 274350
rect 381338 274294 381408 274350
rect 381088 274226 381408 274294
rect 381088 274170 381158 274226
rect 381214 274170 381282 274226
rect 381338 274170 381408 274226
rect 381088 274102 381408 274170
rect 381088 274046 381158 274102
rect 381214 274046 381282 274102
rect 381338 274046 381408 274102
rect 381088 273978 381408 274046
rect 381088 273922 381158 273978
rect 381214 273922 381282 273978
rect 381338 273922 381408 273978
rect 381088 273888 381408 273922
rect 411808 274350 412128 274384
rect 411808 274294 411878 274350
rect 411934 274294 412002 274350
rect 412058 274294 412128 274350
rect 411808 274226 412128 274294
rect 411808 274170 411878 274226
rect 411934 274170 412002 274226
rect 412058 274170 412128 274226
rect 411808 274102 412128 274170
rect 411808 274046 411878 274102
rect 411934 274046 412002 274102
rect 412058 274046 412128 274102
rect 411808 273978 412128 274046
rect 411808 273922 411878 273978
rect 411934 273922 412002 273978
rect 412058 273922 412128 273978
rect 411808 273888 412128 273922
rect 442528 274350 442848 274384
rect 442528 274294 442598 274350
rect 442654 274294 442722 274350
rect 442778 274294 442848 274350
rect 442528 274226 442848 274294
rect 442528 274170 442598 274226
rect 442654 274170 442722 274226
rect 442778 274170 442848 274226
rect 442528 274102 442848 274170
rect 442528 274046 442598 274102
rect 442654 274046 442722 274102
rect 442778 274046 442848 274102
rect 442528 273978 442848 274046
rect 442528 273922 442598 273978
rect 442654 273922 442722 273978
rect 442778 273922 442848 273978
rect 442528 273888 442848 273922
rect 473248 274350 473568 274384
rect 473248 274294 473318 274350
rect 473374 274294 473442 274350
rect 473498 274294 473568 274350
rect 473248 274226 473568 274294
rect 473248 274170 473318 274226
rect 473374 274170 473442 274226
rect 473498 274170 473568 274226
rect 473248 274102 473568 274170
rect 473248 274046 473318 274102
rect 473374 274046 473442 274102
rect 473498 274046 473568 274102
rect 473248 273978 473568 274046
rect 473248 273922 473318 273978
rect 473374 273922 473442 273978
rect 473498 273922 473568 273978
rect 473248 273888 473568 273922
rect 503968 274350 504288 274384
rect 503968 274294 504038 274350
rect 504094 274294 504162 274350
rect 504218 274294 504288 274350
rect 503968 274226 504288 274294
rect 503968 274170 504038 274226
rect 504094 274170 504162 274226
rect 504218 274170 504288 274226
rect 503968 274102 504288 274170
rect 503968 274046 504038 274102
rect 504094 274046 504162 274102
rect 504218 274046 504288 274102
rect 503968 273978 504288 274046
rect 503968 273922 504038 273978
rect 504094 273922 504162 273978
rect 504218 273922 504288 273978
rect 503968 273888 504288 273922
rect 534688 274350 535008 274384
rect 534688 274294 534758 274350
rect 534814 274294 534882 274350
rect 534938 274294 535008 274350
rect 534688 274226 535008 274294
rect 534688 274170 534758 274226
rect 534814 274170 534882 274226
rect 534938 274170 535008 274226
rect 534688 274102 535008 274170
rect 534688 274046 534758 274102
rect 534814 274046 534882 274102
rect 534938 274046 535008 274102
rect 534688 273978 535008 274046
rect 534688 273922 534758 273978
rect 534814 273922 534882 273978
rect 534938 273922 535008 273978
rect 534688 273888 535008 273922
rect 565408 274350 565728 274384
rect 565408 274294 565478 274350
rect 565534 274294 565602 274350
rect 565658 274294 565728 274350
rect 565408 274226 565728 274294
rect 565408 274170 565478 274226
rect 565534 274170 565602 274226
rect 565658 274170 565728 274226
rect 565408 274102 565728 274170
rect 565408 274046 565478 274102
rect 565534 274046 565602 274102
rect 565658 274046 565728 274102
rect 565408 273978 565728 274046
rect 565408 273922 565478 273978
rect 565534 273922 565602 273978
rect 565658 273922 565728 273978
rect 565408 273888 565728 273922
rect 585452 271460 585508 271470
rect 5418 256294 5514 256350
rect 5570 256294 5638 256350
rect 5694 256294 5762 256350
rect 5818 256294 5886 256350
rect 5942 256294 6038 256350
rect 5418 256226 6038 256294
rect 5418 256170 5514 256226
rect 5570 256170 5638 256226
rect 5694 256170 5762 256226
rect 5818 256170 5886 256226
rect 5942 256170 6038 256226
rect 5418 256102 6038 256170
rect 5418 256046 5514 256102
rect 5570 256046 5638 256102
rect 5694 256046 5762 256102
rect 5818 256046 5886 256102
rect 5942 256046 6038 256102
rect 5418 255978 6038 256046
rect 5418 255922 5514 255978
rect 5570 255922 5638 255978
rect 5694 255922 5762 255978
rect 5818 255922 5886 255978
rect 5942 255922 6038 255978
rect 5418 238350 6038 255922
rect 6188 262612 6244 262622
rect 6188 249284 6244 262556
rect 27808 262350 28128 262384
rect 27808 262294 27878 262350
rect 27934 262294 28002 262350
rect 28058 262294 28128 262350
rect 27808 262226 28128 262294
rect 27808 262170 27878 262226
rect 27934 262170 28002 262226
rect 28058 262170 28128 262226
rect 27808 262102 28128 262170
rect 27808 262046 27878 262102
rect 27934 262046 28002 262102
rect 28058 262046 28128 262102
rect 27808 261978 28128 262046
rect 27808 261922 27878 261978
rect 27934 261922 28002 261978
rect 28058 261922 28128 261978
rect 27808 261888 28128 261922
rect 58528 262350 58848 262384
rect 58528 262294 58598 262350
rect 58654 262294 58722 262350
rect 58778 262294 58848 262350
rect 58528 262226 58848 262294
rect 58528 262170 58598 262226
rect 58654 262170 58722 262226
rect 58778 262170 58848 262226
rect 58528 262102 58848 262170
rect 58528 262046 58598 262102
rect 58654 262046 58722 262102
rect 58778 262046 58848 262102
rect 58528 261978 58848 262046
rect 58528 261922 58598 261978
rect 58654 261922 58722 261978
rect 58778 261922 58848 261978
rect 58528 261888 58848 261922
rect 89248 262350 89568 262384
rect 89248 262294 89318 262350
rect 89374 262294 89442 262350
rect 89498 262294 89568 262350
rect 89248 262226 89568 262294
rect 89248 262170 89318 262226
rect 89374 262170 89442 262226
rect 89498 262170 89568 262226
rect 89248 262102 89568 262170
rect 89248 262046 89318 262102
rect 89374 262046 89442 262102
rect 89498 262046 89568 262102
rect 89248 261978 89568 262046
rect 89248 261922 89318 261978
rect 89374 261922 89442 261978
rect 89498 261922 89568 261978
rect 89248 261888 89568 261922
rect 119968 262350 120288 262384
rect 119968 262294 120038 262350
rect 120094 262294 120162 262350
rect 120218 262294 120288 262350
rect 119968 262226 120288 262294
rect 119968 262170 120038 262226
rect 120094 262170 120162 262226
rect 120218 262170 120288 262226
rect 119968 262102 120288 262170
rect 119968 262046 120038 262102
rect 120094 262046 120162 262102
rect 120218 262046 120288 262102
rect 119968 261978 120288 262046
rect 119968 261922 120038 261978
rect 120094 261922 120162 261978
rect 120218 261922 120288 261978
rect 119968 261888 120288 261922
rect 150688 262350 151008 262384
rect 150688 262294 150758 262350
rect 150814 262294 150882 262350
rect 150938 262294 151008 262350
rect 150688 262226 151008 262294
rect 150688 262170 150758 262226
rect 150814 262170 150882 262226
rect 150938 262170 151008 262226
rect 150688 262102 151008 262170
rect 150688 262046 150758 262102
rect 150814 262046 150882 262102
rect 150938 262046 151008 262102
rect 150688 261978 151008 262046
rect 150688 261922 150758 261978
rect 150814 261922 150882 261978
rect 150938 261922 151008 261978
rect 150688 261888 151008 261922
rect 181408 262350 181728 262384
rect 181408 262294 181478 262350
rect 181534 262294 181602 262350
rect 181658 262294 181728 262350
rect 181408 262226 181728 262294
rect 181408 262170 181478 262226
rect 181534 262170 181602 262226
rect 181658 262170 181728 262226
rect 181408 262102 181728 262170
rect 181408 262046 181478 262102
rect 181534 262046 181602 262102
rect 181658 262046 181728 262102
rect 181408 261978 181728 262046
rect 181408 261922 181478 261978
rect 181534 261922 181602 261978
rect 181658 261922 181728 261978
rect 181408 261888 181728 261922
rect 212128 262350 212448 262384
rect 212128 262294 212198 262350
rect 212254 262294 212322 262350
rect 212378 262294 212448 262350
rect 212128 262226 212448 262294
rect 212128 262170 212198 262226
rect 212254 262170 212322 262226
rect 212378 262170 212448 262226
rect 212128 262102 212448 262170
rect 212128 262046 212198 262102
rect 212254 262046 212322 262102
rect 212378 262046 212448 262102
rect 212128 261978 212448 262046
rect 212128 261922 212198 261978
rect 212254 261922 212322 261978
rect 212378 261922 212448 261978
rect 212128 261888 212448 261922
rect 242848 262350 243168 262384
rect 242848 262294 242918 262350
rect 242974 262294 243042 262350
rect 243098 262294 243168 262350
rect 242848 262226 243168 262294
rect 242848 262170 242918 262226
rect 242974 262170 243042 262226
rect 243098 262170 243168 262226
rect 242848 262102 243168 262170
rect 242848 262046 242918 262102
rect 242974 262046 243042 262102
rect 243098 262046 243168 262102
rect 242848 261978 243168 262046
rect 242848 261922 242918 261978
rect 242974 261922 243042 261978
rect 243098 261922 243168 261978
rect 242848 261888 243168 261922
rect 273568 262350 273888 262384
rect 273568 262294 273638 262350
rect 273694 262294 273762 262350
rect 273818 262294 273888 262350
rect 273568 262226 273888 262294
rect 273568 262170 273638 262226
rect 273694 262170 273762 262226
rect 273818 262170 273888 262226
rect 273568 262102 273888 262170
rect 273568 262046 273638 262102
rect 273694 262046 273762 262102
rect 273818 262046 273888 262102
rect 273568 261978 273888 262046
rect 273568 261922 273638 261978
rect 273694 261922 273762 261978
rect 273818 261922 273888 261978
rect 273568 261888 273888 261922
rect 304288 262350 304608 262384
rect 304288 262294 304358 262350
rect 304414 262294 304482 262350
rect 304538 262294 304608 262350
rect 304288 262226 304608 262294
rect 304288 262170 304358 262226
rect 304414 262170 304482 262226
rect 304538 262170 304608 262226
rect 304288 262102 304608 262170
rect 304288 262046 304358 262102
rect 304414 262046 304482 262102
rect 304538 262046 304608 262102
rect 304288 261978 304608 262046
rect 304288 261922 304358 261978
rect 304414 261922 304482 261978
rect 304538 261922 304608 261978
rect 304288 261888 304608 261922
rect 335008 262350 335328 262384
rect 335008 262294 335078 262350
rect 335134 262294 335202 262350
rect 335258 262294 335328 262350
rect 335008 262226 335328 262294
rect 335008 262170 335078 262226
rect 335134 262170 335202 262226
rect 335258 262170 335328 262226
rect 335008 262102 335328 262170
rect 335008 262046 335078 262102
rect 335134 262046 335202 262102
rect 335258 262046 335328 262102
rect 335008 261978 335328 262046
rect 335008 261922 335078 261978
rect 335134 261922 335202 261978
rect 335258 261922 335328 261978
rect 335008 261888 335328 261922
rect 365728 262350 366048 262384
rect 365728 262294 365798 262350
rect 365854 262294 365922 262350
rect 365978 262294 366048 262350
rect 365728 262226 366048 262294
rect 365728 262170 365798 262226
rect 365854 262170 365922 262226
rect 365978 262170 366048 262226
rect 365728 262102 366048 262170
rect 365728 262046 365798 262102
rect 365854 262046 365922 262102
rect 365978 262046 366048 262102
rect 365728 261978 366048 262046
rect 365728 261922 365798 261978
rect 365854 261922 365922 261978
rect 365978 261922 366048 261978
rect 365728 261888 366048 261922
rect 396448 262350 396768 262384
rect 396448 262294 396518 262350
rect 396574 262294 396642 262350
rect 396698 262294 396768 262350
rect 396448 262226 396768 262294
rect 396448 262170 396518 262226
rect 396574 262170 396642 262226
rect 396698 262170 396768 262226
rect 396448 262102 396768 262170
rect 396448 262046 396518 262102
rect 396574 262046 396642 262102
rect 396698 262046 396768 262102
rect 396448 261978 396768 262046
rect 396448 261922 396518 261978
rect 396574 261922 396642 261978
rect 396698 261922 396768 261978
rect 396448 261888 396768 261922
rect 427168 262350 427488 262384
rect 427168 262294 427238 262350
rect 427294 262294 427362 262350
rect 427418 262294 427488 262350
rect 427168 262226 427488 262294
rect 427168 262170 427238 262226
rect 427294 262170 427362 262226
rect 427418 262170 427488 262226
rect 427168 262102 427488 262170
rect 427168 262046 427238 262102
rect 427294 262046 427362 262102
rect 427418 262046 427488 262102
rect 427168 261978 427488 262046
rect 427168 261922 427238 261978
rect 427294 261922 427362 261978
rect 427418 261922 427488 261978
rect 427168 261888 427488 261922
rect 457888 262350 458208 262384
rect 457888 262294 457958 262350
rect 458014 262294 458082 262350
rect 458138 262294 458208 262350
rect 457888 262226 458208 262294
rect 457888 262170 457958 262226
rect 458014 262170 458082 262226
rect 458138 262170 458208 262226
rect 457888 262102 458208 262170
rect 457888 262046 457958 262102
rect 458014 262046 458082 262102
rect 458138 262046 458208 262102
rect 457888 261978 458208 262046
rect 457888 261922 457958 261978
rect 458014 261922 458082 261978
rect 458138 261922 458208 261978
rect 457888 261888 458208 261922
rect 488608 262350 488928 262384
rect 488608 262294 488678 262350
rect 488734 262294 488802 262350
rect 488858 262294 488928 262350
rect 488608 262226 488928 262294
rect 488608 262170 488678 262226
rect 488734 262170 488802 262226
rect 488858 262170 488928 262226
rect 488608 262102 488928 262170
rect 488608 262046 488678 262102
rect 488734 262046 488802 262102
rect 488858 262046 488928 262102
rect 488608 261978 488928 262046
rect 488608 261922 488678 261978
rect 488734 261922 488802 261978
rect 488858 261922 488928 261978
rect 488608 261888 488928 261922
rect 519328 262350 519648 262384
rect 519328 262294 519398 262350
rect 519454 262294 519522 262350
rect 519578 262294 519648 262350
rect 519328 262226 519648 262294
rect 519328 262170 519398 262226
rect 519454 262170 519522 262226
rect 519578 262170 519648 262226
rect 519328 262102 519648 262170
rect 519328 262046 519398 262102
rect 519454 262046 519522 262102
rect 519578 262046 519648 262102
rect 519328 261978 519648 262046
rect 519328 261922 519398 261978
rect 519454 261922 519522 261978
rect 519578 261922 519648 261978
rect 519328 261888 519648 261922
rect 550048 262350 550368 262384
rect 550048 262294 550118 262350
rect 550174 262294 550242 262350
rect 550298 262294 550368 262350
rect 550048 262226 550368 262294
rect 550048 262170 550118 262226
rect 550174 262170 550242 262226
rect 550298 262170 550368 262226
rect 550048 262102 550368 262170
rect 550048 262046 550118 262102
rect 550174 262046 550242 262102
rect 550298 262046 550368 262102
rect 550048 261978 550368 262046
rect 550048 261922 550118 261978
rect 550174 261922 550242 261978
rect 550298 261922 550368 261978
rect 550048 261888 550368 261922
rect 12448 256350 12768 256384
rect 12448 256294 12518 256350
rect 12574 256294 12642 256350
rect 12698 256294 12768 256350
rect 12448 256226 12768 256294
rect 12448 256170 12518 256226
rect 12574 256170 12642 256226
rect 12698 256170 12768 256226
rect 12448 256102 12768 256170
rect 12448 256046 12518 256102
rect 12574 256046 12642 256102
rect 12698 256046 12768 256102
rect 12448 255978 12768 256046
rect 12448 255922 12518 255978
rect 12574 255922 12642 255978
rect 12698 255922 12768 255978
rect 12448 255888 12768 255922
rect 43168 256350 43488 256384
rect 43168 256294 43238 256350
rect 43294 256294 43362 256350
rect 43418 256294 43488 256350
rect 43168 256226 43488 256294
rect 43168 256170 43238 256226
rect 43294 256170 43362 256226
rect 43418 256170 43488 256226
rect 43168 256102 43488 256170
rect 43168 256046 43238 256102
rect 43294 256046 43362 256102
rect 43418 256046 43488 256102
rect 43168 255978 43488 256046
rect 43168 255922 43238 255978
rect 43294 255922 43362 255978
rect 43418 255922 43488 255978
rect 43168 255888 43488 255922
rect 73888 256350 74208 256384
rect 73888 256294 73958 256350
rect 74014 256294 74082 256350
rect 74138 256294 74208 256350
rect 73888 256226 74208 256294
rect 73888 256170 73958 256226
rect 74014 256170 74082 256226
rect 74138 256170 74208 256226
rect 73888 256102 74208 256170
rect 73888 256046 73958 256102
rect 74014 256046 74082 256102
rect 74138 256046 74208 256102
rect 73888 255978 74208 256046
rect 73888 255922 73958 255978
rect 74014 255922 74082 255978
rect 74138 255922 74208 255978
rect 73888 255888 74208 255922
rect 104608 256350 104928 256384
rect 104608 256294 104678 256350
rect 104734 256294 104802 256350
rect 104858 256294 104928 256350
rect 104608 256226 104928 256294
rect 104608 256170 104678 256226
rect 104734 256170 104802 256226
rect 104858 256170 104928 256226
rect 104608 256102 104928 256170
rect 104608 256046 104678 256102
rect 104734 256046 104802 256102
rect 104858 256046 104928 256102
rect 104608 255978 104928 256046
rect 104608 255922 104678 255978
rect 104734 255922 104802 255978
rect 104858 255922 104928 255978
rect 104608 255888 104928 255922
rect 135328 256350 135648 256384
rect 135328 256294 135398 256350
rect 135454 256294 135522 256350
rect 135578 256294 135648 256350
rect 135328 256226 135648 256294
rect 135328 256170 135398 256226
rect 135454 256170 135522 256226
rect 135578 256170 135648 256226
rect 135328 256102 135648 256170
rect 135328 256046 135398 256102
rect 135454 256046 135522 256102
rect 135578 256046 135648 256102
rect 135328 255978 135648 256046
rect 135328 255922 135398 255978
rect 135454 255922 135522 255978
rect 135578 255922 135648 255978
rect 135328 255888 135648 255922
rect 166048 256350 166368 256384
rect 166048 256294 166118 256350
rect 166174 256294 166242 256350
rect 166298 256294 166368 256350
rect 166048 256226 166368 256294
rect 166048 256170 166118 256226
rect 166174 256170 166242 256226
rect 166298 256170 166368 256226
rect 166048 256102 166368 256170
rect 166048 256046 166118 256102
rect 166174 256046 166242 256102
rect 166298 256046 166368 256102
rect 166048 255978 166368 256046
rect 166048 255922 166118 255978
rect 166174 255922 166242 255978
rect 166298 255922 166368 255978
rect 166048 255888 166368 255922
rect 196768 256350 197088 256384
rect 196768 256294 196838 256350
rect 196894 256294 196962 256350
rect 197018 256294 197088 256350
rect 196768 256226 197088 256294
rect 196768 256170 196838 256226
rect 196894 256170 196962 256226
rect 197018 256170 197088 256226
rect 196768 256102 197088 256170
rect 196768 256046 196838 256102
rect 196894 256046 196962 256102
rect 197018 256046 197088 256102
rect 196768 255978 197088 256046
rect 196768 255922 196838 255978
rect 196894 255922 196962 255978
rect 197018 255922 197088 255978
rect 196768 255888 197088 255922
rect 227488 256350 227808 256384
rect 227488 256294 227558 256350
rect 227614 256294 227682 256350
rect 227738 256294 227808 256350
rect 227488 256226 227808 256294
rect 227488 256170 227558 256226
rect 227614 256170 227682 256226
rect 227738 256170 227808 256226
rect 227488 256102 227808 256170
rect 227488 256046 227558 256102
rect 227614 256046 227682 256102
rect 227738 256046 227808 256102
rect 227488 255978 227808 256046
rect 227488 255922 227558 255978
rect 227614 255922 227682 255978
rect 227738 255922 227808 255978
rect 227488 255888 227808 255922
rect 258208 256350 258528 256384
rect 258208 256294 258278 256350
rect 258334 256294 258402 256350
rect 258458 256294 258528 256350
rect 258208 256226 258528 256294
rect 258208 256170 258278 256226
rect 258334 256170 258402 256226
rect 258458 256170 258528 256226
rect 258208 256102 258528 256170
rect 258208 256046 258278 256102
rect 258334 256046 258402 256102
rect 258458 256046 258528 256102
rect 258208 255978 258528 256046
rect 258208 255922 258278 255978
rect 258334 255922 258402 255978
rect 258458 255922 258528 255978
rect 258208 255888 258528 255922
rect 288928 256350 289248 256384
rect 288928 256294 288998 256350
rect 289054 256294 289122 256350
rect 289178 256294 289248 256350
rect 288928 256226 289248 256294
rect 288928 256170 288998 256226
rect 289054 256170 289122 256226
rect 289178 256170 289248 256226
rect 288928 256102 289248 256170
rect 288928 256046 288998 256102
rect 289054 256046 289122 256102
rect 289178 256046 289248 256102
rect 288928 255978 289248 256046
rect 288928 255922 288998 255978
rect 289054 255922 289122 255978
rect 289178 255922 289248 255978
rect 288928 255888 289248 255922
rect 319648 256350 319968 256384
rect 319648 256294 319718 256350
rect 319774 256294 319842 256350
rect 319898 256294 319968 256350
rect 319648 256226 319968 256294
rect 319648 256170 319718 256226
rect 319774 256170 319842 256226
rect 319898 256170 319968 256226
rect 319648 256102 319968 256170
rect 319648 256046 319718 256102
rect 319774 256046 319842 256102
rect 319898 256046 319968 256102
rect 319648 255978 319968 256046
rect 319648 255922 319718 255978
rect 319774 255922 319842 255978
rect 319898 255922 319968 255978
rect 319648 255888 319968 255922
rect 350368 256350 350688 256384
rect 350368 256294 350438 256350
rect 350494 256294 350562 256350
rect 350618 256294 350688 256350
rect 350368 256226 350688 256294
rect 350368 256170 350438 256226
rect 350494 256170 350562 256226
rect 350618 256170 350688 256226
rect 350368 256102 350688 256170
rect 350368 256046 350438 256102
rect 350494 256046 350562 256102
rect 350618 256046 350688 256102
rect 350368 255978 350688 256046
rect 350368 255922 350438 255978
rect 350494 255922 350562 255978
rect 350618 255922 350688 255978
rect 350368 255888 350688 255922
rect 381088 256350 381408 256384
rect 381088 256294 381158 256350
rect 381214 256294 381282 256350
rect 381338 256294 381408 256350
rect 381088 256226 381408 256294
rect 381088 256170 381158 256226
rect 381214 256170 381282 256226
rect 381338 256170 381408 256226
rect 381088 256102 381408 256170
rect 381088 256046 381158 256102
rect 381214 256046 381282 256102
rect 381338 256046 381408 256102
rect 381088 255978 381408 256046
rect 381088 255922 381158 255978
rect 381214 255922 381282 255978
rect 381338 255922 381408 255978
rect 381088 255888 381408 255922
rect 411808 256350 412128 256384
rect 411808 256294 411878 256350
rect 411934 256294 412002 256350
rect 412058 256294 412128 256350
rect 411808 256226 412128 256294
rect 411808 256170 411878 256226
rect 411934 256170 412002 256226
rect 412058 256170 412128 256226
rect 411808 256102 412128 256170
rect 411808 256046 411878 256102
rect 411934 256046 412002 256102
rect 412058 256046 412128 256102
rect 411808 255978 412128 256046
rect 411808 255922 411878 255978
rect 411934 255922 412002 255978
rect 412058 255922 412128 255978
rect 411808 255888 412128 255922
rect 442528 256350 442848 256384
rect 442528 256294 442598 256350
rect 442654 256294 442722 256350
rect 442778 256294 442848 256350
rect 442528 256226 442848 256294
rect 442528 256170 442598 256226
rect 442654 256170 442722 256226
rect 442778 256170 442848 256226
rect 442528 256102 442848 256170
rect 442528 256046 442598 256102
rect 442654 256046 442722 256102
rect 442778 256046 442848 256102
rect 442528 255978 442848 256046
rect 442528 255922 442598 255978
rect 442654 255922 442722 255978
rect 442778 255922 442848 255978
rect 442528 255888 442848 255922
rect 473248 256350 473568 256384
rect 473248 256294 473318 256350
rect 473374 256294 473442 256350
rect 473498 256294 473568 256350
rect 473248 256226 473568 256294
rect 473248 256170 473318 256226
rect 473374 256170 473442 256226
rect 473498 256170 473568 256226
rect 473248 256102 473568 256170
rect 473248 256046 473318 256102
rect 473374 256046 473442 256102
rect 473498 256046 473568 256102
rect 473248 255978 473568 256046
rect 473248 255922 473318 255978
rect 473374 255922 473442 255978
rect 473498 255922 473568 255978
rect 473248 255888 473568 255922
rect 503968 256350 504288 256384
rect 503968 256294 504038 256350
rect 504094 256294 504162 256350
rect 504218 256294 504288 256350
rect 503968 256226 504288 256294
rect 503968 256170 504038 256226
rect 504094 256170 504162 256226
rect 504218 256170 504288 256226
rect 503968 256102 504288 256170
rect 503968 256046 504038 256102
rect 504094 256046 504162 256102
rect 504218 256046 504288 256102
rect 503968 255978 504288 256046
rect 503968 255922 504038 255978
rect 504094 255922 504162 255978
rect 504218 255922 504288 255978
rect 503968 255888 504288 255922
rect 534688 256350 535008 256384
rect 534688 256294 534758 256350
rect 534814 256294 534882 256350
rect 534938 256294 535008 256350
rect 534688 256226 535008 256294
rect 534688 256170 534758 256226
rect 534814 256170 534882 256226
rect 534938 256170 535008 256226
rect 534688 256102 535008 256170
rect 534688 256046 534758 256102
rect 534814 256046 534882 256102
rect 534938 256046 535008 256102
rect 534688 255978 535008 256046
rect 534688 255922 534758 255978
rect 534814 255922 534882 255978
rect 534938 255922 535008 255978
rect 534688 255888 535008 255922
rect 565408 256350 565728 256384
rect 565408 256294 565478 256350
rect 565534 256294 565602 256350
rect 565658 256294 565728 256350
rect 565408 256226 565728 256294
rect 565408 256170 565478 256226
rect 565534 256170 565602 256226
rect 565658 256170 565728 256226
rect 565408 256102 565728 256170
rect 565408 256046 565478 256102
rect 565534 256046 565602 256102
rect 565658 256046 565728 256102
rect 565408 255978 565728 256046
rect 565408 255922 565478 255978
rect 565534 255922 565602 255978
rect 565658 255922 565728 255978
rect 565408 255888 565728 255922
rect 6188 249218 6244 249228
rect 5418 238294 5514 238350
rect 5570 238294 5638 238350
rect 5694 238294 5762 238350
rect 5818 238294 5886 238350
rect 5942 238294 6038 238350
rect 5418 238226 6038 238294
rect 5418 238170 5514 238226
rect 5570 238170 5638 238226
rect 5694 238170 5762 238226
rect 5818 238170 5886 238226
rect 5942 238170 6038 238226
rect 5418 238102 6038 238170
rect 5418 238046 5514 238102
rect 5570 238046 5638 238102
rect 5694 238046 5762 238102
rect 5818 238046 5886 238102
rect 5942 238046 6038 238102
rect 5418 237978 6038 238046
rect 5418 237922 5514 237978
rect 5570 237922 5638 237978
rect 5694 237922 5762 237978
rect 5818 237922 5886 237978
rect 5942 237922 6038 237978
rect -956 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 -336 220350
rect -956 220226 -336 220294
rect -956 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 -336 220226
rect -956 220102 -336 220170
rect -956 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 -336 220102
rect -956 219978 -336 220046
rect -956 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 -336 219978
rect -956 202350 -336 219922
rect 4172 234388 4228 234398
rect 4172 217700 4228 234332
rect 4172 217634 4228 217644
rect 5418 220350 6038 237922
rect 6188 248500 6244 248510
rect 6188 228228 6244 248444
rect 27808 244350 28128 244384
rect 27808 244294 27878 244350
rect 27934 244294 28002 244350
rect 28058 244294 28128 244350
rect 27808 244226 28128 244294
rect 27808 244170 27878 244226
rect 27934 244170 28002 244226
rect 28058 244170 28128 244226
rect 27808 244102 28128 244170
rect 27808 244046 27878 244102
rect 27934 244046 28002 244102
rect 28058 244046 28128 244102
rect 27808 243978 28128 244046
rect 27808 243922 27878 243978
rect 27934 243922 28002 243978
rect 28058 243922 28128 243978
rect 27808 243888 28128 243922
rect 58528 244350 58848 244384
rect 58528 244294 58598 244350
rect 58654 244294 58722 244350
rect 58778 244294 58848 244350
rect 58528 244226 58848 244294
rect 58528 244170 58598 244226
rect 58654 244170 58722 244226
rect 58778 244170 58848 244226
rect 58528 244102 58848 244170
rect 58528 244046 58598 244102
rect 58654 244046 58722 244102
rect 58778 244046 58848 244102
rect 58528 243978 58848 244046
rect 58528 243922 58598 243978
rect 58654 243922 58722 243978
rect 58778 243922 58848 243978
rect 58528 243888 58848 243922
rect 89248 244350 89568 244384
rect 89248 244294 89318 244350
rect 89374 244294 89442 244350
rect 89498 244294 89568 244350
rect 89248 244226 89568 244294
rect 89248 244170 89318 244226
rect 89374 244170 89442 244226
rect 89498 244170 89568 244226
rect 89248 244102 89568 244170
rect 89248 244046 89318 244102
rect 89374 244046 89442 244102
rect 89498 244046 89568 244102
rect 89248 243978 89568 244046
rect 89248 243922 89318 243978
rect 89374 243922 89442 243978
rect 89498 243922 89568 243978
rect 89248 243888 89568 243922
rect 119968 244350 120288 244384
rect 119968 244294 120038 244350
rect 120094 244294 120162 244350
rect 120218 244294 120288 244350
rect 119968 244226 120288 244294
rect 119968 244170 120038 244226
rect 120094 244170 120162 244226
rect 120218 244170 120288 244226
rect 119968 244102 120288 244170
rect 119968 244046 120038 244102
rect 120094 244046 120162 244102
rect 120218 244046 120288 244102
rect 119968 243978 120288 244046
rect 119968 243922 120038 243978
rect 120094 243922 120162 243978
rect 120218 243922 120288 243978
rect 119968 243888 120288 243922
rect 150688 244350 151008 244384
rect 150688 244294 150758 244350
rect 150814 244294 150882 244350
rect 150938 244294 151008 244350
rect 150688 244226 151008 244294
rect 150688 244170 150758 244226
rect 150814 244170 150882 244226
rect 150938 244170 151008 244226
rect 150688 244102 151008 244170
rect 150688 244046 150758 244102
rect 150814 244046 150882 244102
rect 150938 244046 151008 244102
rect 150688 243978 151008 244046
rect 150688 243922 150758 243978
rect 150814 243922 150882 243978
rect 150938 243922 151008 243978
rect 150688 243888 151008 243922
rect 181408 244350 181728 244384
rect 181408 244294 181478 244350
rect 181534 244294 181602 244350
rect 181658 244294 181728 244350
rect 181408 244226 181728 244294
rect 181408 244170 181478 244226
rect 181534 244170 181602 244226
rect 181658 244170 181728 244226
rect 181408 244102 181728 244170
rect 181408 244046 181478 244102
rect 181534 244046 181602 244102
rect 181658 244046 181728 244102
rect 181408 243978 181728 244046
rect 181408 243922 181478 243978
rect 181534 243922 181602 243978
rect 181658 243922 181728 243978
rect 181408 243888 181728 243922
rect 212128 244350 212448 244384
rect 212128 244294 212198 244350
rect 212254 244294 212322 244350
rect 212378 244294 212448 244350
rect 212128 244226 212448 244294
rect 212128 244170 212198 244226
rect 212254 244170 212322 244226
rect 212378 244170 212448 244226
rect 212128 244102 212448 244170
rect 212128 244046 212198 244102
rect 212254 244046 212322 244102
rect 212378 244046 212448 244102
rect 212128 243978 212448 244046
rect 212128 243922 212198 243978
rect 212254 243922 212322 243978
rect 212378 243922 212448 243978
rect 212128 243888 212448 243922
rect 242848 244350 243168 244384
rect 242848 244294 242918 244350
rect 242974 244294 243042 244350
rect 243098 244294 243168 244350
rect 242848 244226 243168 244294
rect 242848 244170 242918 244226
rect 242974 244170 243042 244226
rect 243098 244170 243168 244226
rect 242848 244102 243168 244170
rect 242848 244046 242918 244102
rect 242974 244046 243042 244102
rect 243098 244046 243168 244102
rect 242848 243978 243168 244046
rect 242848 243922 242918 243978
rect 242974 243922 243042 243978
rect 243098 243922 243168 243978
rect 242848 243888 243168 243922
rect 273568 244350 273888 244384
rect 273568 244294 273638 244350
rect 273694 244294 273762 244350
rect 273818 244294 273888 244350
rect 273568 244226 273888 244294
rect 273568 244170 273638 244226
rect 273694 244170 273762 244226
rect 273818 244170 273888 244226
rect 273568 244102 273888 244170
rect 273568 244046 273638 244102
rect 273694 244046 273762 244102
rect 273818 244046 273888 244102
rect 273568 243978 273888 244046
rect 273568 243922 273638 243978
rect 273694 243922 273762 243978
rect 273818 243922 273888 243978
rect 273568 243888 273888 243922
rect 304288 244350 304608 244384
rect 304288 244294 304358 244350
rect 304414 244294 304482 244350
rect 304538 244294 304608 244350
rect 304288 244226 304608 244294
rect 304288 244170 304358 244226
rect 304414 244170 304482 244226
rect 304538 244170 304608 244226
rect 304288 244102 304608 244170
rect 304288 244046 304358 244102
rect 304414 244046 304482 244102
rect 304538 244046 304608 244102
rect 304288 243978 304608 244046
rect 304288 243922 304358 243978
rect 304414 243922 304482 243978
rect 304538 243922 304608 243978
rect 304288 243888 304608 243922
rect 335008 244350 335328 244384
rect 335008 244294 335078 244350
rect 335134 244294 335202 244350
rect 335258 244294 335328 244350
rect 335008 244226 335328 244294
rect 335008 244170 335078 244226
rect 335134 244170 335202 244226
rect 335258 244170 335328 244226
rect 335008 244102 335328 244170
rect 335008 244046 335078 244102
rect 335134 244046 335202 244102
rect 335258 244046 335328 244102
rect 335008 243978 335328 244046
rect 335008 243922 335078 243978
rect 335134 243922 335202 243978
rect 335258 243922 335328 243978
rect 335008 243888 335328 243922
rect 365728 244350 366048 244384
rect 365728 244294 365798 244350
rect 365854 244294 365922 244350
rect 365978 244294 366048 244350
rect 365728 244226 366048 244294
rect 365728 244170 365798 244226
rect 365854 244170 365922 244226
rect 365978 244170 366048 244226
rect 365728 244102 366048 244170
rect 365728 244046 365798 244102
rect 365854 244046 365922 244102
rect 365978 244046 366048 244102
rect 365728 243978 366048 244046
rect 365728 243922 365798 243978
rect 365854 243922 365922 243978
rect 365978 243922 366048 243978
rect 365728 243888 366048 243922
rect 396448 244350 396768 244384
rect 396448 244294 396518 244350
rect 396574 244294 396642 244350
rect 396698 244294 396768 244350
rect 396448 244226 396768 244294
rect 396448 244170 396518 244226
rect 396574 244170 396642 244226
rect 396698 244170 396768 244226
rect 396448 244102 396768 244170
rect 396448 244046 396518 244102
rect 396574 244046 396642 244102
rect 396698 244046 396768 244102
rect 396448 243978 396768 244046
rect 396448 243922 396518 243978
rect 396574 243922 396642 243978
rect 396698 243922 396768 243978
rect 396448 243888 396768 243922
rect 427168 244350 427488 244384
rect 427168 244294 427238 244350
rect 427294 244294 427362 244350
rect 427418 244294 427488 244350
rect 427168 244226 427488 244294
rect 427168 244170 427238 244226
rect 427294 244170 427362 244226
rect 427418 244170 427488 244226
rect 427168 244102 427488 244170
rect 427168 244046 427238 244102
rect 427294 244046 427362 244102
rect 427418 244046 427488 244102
rect 427168 243978 427488 244046
rect 427168 243922 427238 243978
rect 427294 243922 427362 243978
rect 427418 243922 427488 243978
rect 427168 243888 427488 243922
rect 457888 244350 458208 244384
rect 457888 244294 457958 244350
rect 458014 244294 458082 244350
rect 458138 244294 458208 244350
rect 457888 244226 458208 244294
rect 457888 244170 457958 244226
rect 458014 244170 458082 244226
rect 458138 244170 458208 244226
rect 457888 244102 458208 244170
rect 457888 244046 457958 244102
rect 458014 244046 458082 244102
rect 458138 244046 458208 244102
rect 457888 243978 458208 244046
rect 457888 243922 457958 243978
rect 458014 243922 458082 243978
rect 458138 243922 458208 243978
rect 457888 243888 458208 243922
rect 488608 244350 488928 244384
rect 488608 244294 488678 244350
rect 488734 244294 488802 244350
rect 488858 244294 488928 244350
rect 488608 244226 488928 244294
rect 488608 244170 488678 244226
rect 488734 244170 488802 244226
rect 488858 244170 488928 244226
rect 488608 244102 488928 244170
rect 488608 244046 488678 244102
rect 488734 244046 488802 244102
rect 488858 244046 488928 244102
rect 488608 243978 488928 244046
rect 488608 243922 488678 243978
rect 488734 243922 488802 243978
rect 488858 243922 488928 243978
rect 488608 243888 488928 243922
rect 519328 244350 519648 244384
rect 519328 244294 519398 244350
rect 519454 244294 519522 244350
rect 519578 244294 519648 244350
rect 519328 244226 519648 244294
rect 519328 244170 519398 244226
rect 519454 244170 519522 244226
rect 519578 244170 519648 244226
rect 519328 244102 519648 244170
rect 519328 244046 519398 244102
rect 519454 244046 519522 244102
rect 519578 244046 519648 244102
rect 519328 243978 519648 244046
rect 519328 243922 519398 243978
rect 519454 243922 519522 243978
rect 519578 243922 519648 243978
rect 519328 243888 519648 243922
rect 550048 244350 550368 244384
rect 550048 244294 550118 244350
rect 550174 244294 550242 244350
rect 550298 244294 550368 244350
rect 550048 244226 550368 244294
rect 550048 244170 550118 244226
rect 550174 244170 550242 244226
rect 550298 244170 550368 244226
rect 550048 244102 550368 244170
rect 550048 244046 550118 244102
rect 550174 244046 550242 244102
rect 550298 244046 550368 244102
rect 550048 243978 550368 244046
rect 550048 243922 550118 243978
rect 550174 243922 550242 243978
rect 550298 243922 550368 243978
rect 550048 243888 550368 243922
rect 12448 238350 12768 238384
rect 12448 238294 12518 238350
rect 12574 238294 12642 238350
rect 12698 238294 12768 238350
rect 12448 238226 12768 238294
rect 12448 238170 12518 238226
rect 12574 238170 12642 238226
rect 12698 238170 12768 238226
rect 12448 238102 12768 238170
rect 12448 238046 12518 238102
rect 12574 238046 12642 238102
rect 12698 238046 12768 238102
rect 12448 237978 12768 238046
rect 12448 237922 12518 237978
rect 12574 237922 12642 237978
rect 12698 237922 12768 237978
rect 12448 237888 12768 237922
rect 43168 238350 43488 238384
rect 43168 238294 43238 238350
rect 43294 238294 43362 238350
rect 43418 238294 43488 238350
rect 43168 238226 43488 238294
rect 43168 238170 43238 238226
rect 43294 238170 43362 238226
rect 43418 238170 43488 238226
rect 43168 238102 43488 238170
rect 43168 238046 43238 238102
rect 43294 238046 43362 238102
rect 43418 238046 43488 238102
rect 43168 237978 43488 238046
rect 43168 237922 43238 237978
rect 43294 237922 43362 237978
rect 43418 237922 43488 237978
rect 43168 237888 43488 237922
rect 73888 238350 74208 238384
rect 73888 238294 73958 238350
rect 74014 238294 74082 238350
rect 74138 238294 74208 238350
rect 73888 238226 74208 238294
rect 73888 238170 73958 238226
rect 74014 238170 74082 238226
rect 74138 238170 74208 238226
rect 73888 238102 74208 238170
rect 73888 238046 73958 238102
rect 74014 238046 74082 238102
rect 74138 238046 74208 238102
rect 73888 237978 74208 238046
rect 73888 237922 73958 237978
rect 74014 237922 74082 237978
rect 74138 237922 74208 237978
rect 73888 237888 74208 237922
rect 104608 238350 104928 238384
rect 104608 238294 104678 238350
rect 104734 238294 104802 238350
rect 104858 238294 104928 238350
rect 104608 238226 104928 238294
rect 104608 238170 104678 238226
rect 104734 238170 104802 238226
rect 104858 238170 104928 238226
rect 104608 238102 104928 238170
rect 104608 238046 104678 238102
rect 104734 238046 104802 238102
rect 104858 238046 104928 238102
rect 104608 237978 104928 238046
rect 104608 237922 104678 237978
rect 104734 237922 104802 237978
rect 104858 237922 104928 237978
rect 104608 237888 104928 237922
rect 135328 238350 135648 238384
rect 135328 238294 135398 238350
rect 135454 238294 135522 238350
rect 135578 238294 135648 238350
rect 135328 238226 135648 238294
rect 135328 238170 135398 238226
rect 135454 238170 135522 238226
rect 135578 238170 135648 238226
rect 135328 238102 135648 238170
rect 135328 238046 135398 238102
rect 135454 238046 135522 238102
rect 135578 238046 135648 238102
rect 135328 237978 135648 238046
rect 135328 237922 135398 237978
rect 135454 237922 135522 237978
rect 135578 237922 135648 237978
rect 135328 237888 135648 237922
rect 166048 238350 166368 238384
rect 166048 238294 166118 238350
rect 166174 238294 166242 238350
rect 166298 238294 166368 238350
rect 166048 238226 166368 238294
rect 166048 238170 166118 238226
rect 166174 238170 166242 238226
rect 166298 238170 166368 238226
rect 166048 238102 166368 238170
rect 166048 238046 166118 238102
rect 166174 238046 166242 238102
rect 166298 238046 166368 238102
rect 166048 237978 166368 238046
rect 166048 237922 166118 237978
rect 166174 237922 166242 237978
rect 166298 237922 166368 237978
rect 166048 237888 166368 237922
rect 196768 238350 197088 238384
rect 196768 238294 196838 238350
rect 196894 238294 196962 238350
rect 197018 238294 197088 238350
rect 196768 238226 197088 238294
rect 196768 238170 196838 238226
rect 196894 238170 196962 238226
rect 197018 238170 197088 238226
rect 196768 238102 197088 238170
rect 196768 238046 196838 238102
rect 196894 238046 196962 238102
rect 197018 238046 197088 238102
rect 196768 237978 197088 238046
rect 196768 237922 196838 237978
rect 196894 237922 196962 237978
rect 197018 237922 197088 237978
rect 196768 237888 197088 237922
rect 227488 238350 227808 238384
rect 227488 238294 227558 238350
rect 227614 238294 227682 238350
rect 227738 238294 227808 238350
rect 227488 238226 227808 238294
rect 227488 238170 227558 238226
rect 227614 238170 227682 238226
rect 227738 238170 227808 238226
rect 227488 238102 227808 238170
rect 227488 238046 227558 238102
rect 227614 238046 227682 238102
rect 227738 238046 227808 238102
rect 227488 237978 227808 238046
rect 227488 237922 227558 237978
rect 227614 237922 227682 237978
rect 227738 237922 227808 237978
rect 227488 237888 227808 237922
rect 258208 238350 258528 238384
rect 258208 238294 258278 238350
rect 258334 238294 258402 238350
rect 258458 238294 258528 238350
rect 258208 238226 258528 238294
rect 258208 238170 258278 238226
rect 258334 238170 258402 238226
rect 258458 238170 258528 238226
rect 258208 238102 258528 238170
rect 258208 238046 258278 238102
rect 258334 238046 258402 238102
rect 258458 238046 258528 238102
rect 258208 237978 258528 238046
rect 258208 237922 258278 237978
rect 258334 237922 258402 237978
rect 258458 237922 258528 237978
rect 258208 237888 258528 237922
rect 288928 238350 289248 238384
rect 288928 238294 288998 238350
rect 289054 238294 289122 238350
rect 289178 238294 289248 238350
rect 288928 238226 289248 238294
rect 288928 238170 288998 238226
rect 289054 238170 289122 238226
rect 289178 238170 289248 238226
rect 288928 238102 289248 238170
rect 288928 238046 288998 238102
rect 289054 238046 289122 238102
rect 289178 238046 289248 238102
rect 288928 237978 289248 238046
rect 288928 237922 288998 237978
rect 289054 237922 289122 237978
rect 289178 237922 289248 237978
rect 288928 237888 289248 237922
rect 319648 238350 319968 238384
rect 319648 238294 319718 238350
rect 319774 238294 319842 238350
rect 319898 238294 319968 238350
rect 319648 238226 319968 238294
rect 319648 238170 319718 238226
rect 319774 238170 319842 238226
rect 319898 238170 319968 238226
rect 319648 238102 319968 238170
rect 319648 238046 319718 238102
rect 319774 238046 319842 238102
rect 319898 238046 319968 238102
rect 319648 237978 319968 238046
rect 319648 237922 319718 237978
rect 319774 237922 319842 237978
rect 319898 237922 319968 237978
rect 319648 237888 319968 237922
rect 350368 238350 350688 238384
rect 350368 238294 350438 238350
rect 350494 238294 350562 238350
rect 350618 238294 350688 238350
rect 350368 238226 350688 238294
rect 350368 238170 350438 238226
rect 350494 238170 350562 238226
rect 350618 238170 350688 238226
rect 350368 238102 350688 238170
rect 350368 238046 350438 238102
rect 350494 238046 350562 238102
rect 350618 238046 350688 238102
rect 350368 237978 350688 238046
rect 350368 237922 350438 237978
rect 350494 237922 350562 237978
rect 350618 237922 350688 237978
rect 350368 237888 350688 237922
rect 381088 238350 381408 238384
rect 381088 238294 381158 238350
rect 381214 238294 381282 238350
rect 381338 238294 381408 238350
rect 381088 238226 381408 238294
rect 381088 238170 381158 238226
rect 381214 238170 381282 238226
rect 381338 238170 381408 238226
rect 381088 238102 381408 238170
rect 381088 238046 381158 238102
rect 381214 238046 381282 238102
rect 381338 238046 381408 238102
rect 381088 237978 381408 238046
rect 381088 237922 381158 237978
rect 381214 237922 381282 237978
rect 381338 237922 381408 237978
rect 381088 237888 381408 237922
rect 411808 238350 412128 238384
rect 411808 238294 411878 238350
rect 411934 238294 412002 238350
rect 412058 238294 412128 238350
rect 411808 238226 412128 238294
rect 411808 238170 411878 238226
rect 411934 238170 412002 238226
rect 412058 238170 412128 238226
rect 411808 238102 412128 238170
rect 411808 238046 411878 238102
rect 411934 238046 412002 238102
rect 412058 238046 412128 238102
rect 411808 237978 412128 238046
rect 411808 237922 411878 237978
rect 411934 237922 412002 237978
rect 412058 237922 412128 237978
rect 411808 237888 412128 237922
rect 442528 238350 442848 238384
rect 442528 238294 442598 238350
rect 442654 238294 442722 238350
rect 442778 238294 442848 238350
rect 442528 238226 442848 238294
rect 442528 238170 442598 238226
rect 442654 238170 442722 238226
rect 442778 238170 442848 238226
rect 442528 238102 442848 238170
rect 442528 238046 442598 238102
rect 442654 238046 442722 238102
rect 442778 238046 442848 238102
rect 442528 237978 442848 238046
rect 442528 237922 442598 237978
rect 442654 237922 442722 237978
rect 442778 237922 442848 237978
rect 442528 237888 442848 237922
rect 473248 238350 473568 238384
rect 473248 238294 473318 238350
rect 473374 238294 473442 238350
rect 473498 238294 473568 238350
rect 473248 238226 473568 238294
rect 473248 238170 473318 238226
rect 473374 238170 473442 238226
rect 473498 238170 473568 238226
rect 473248 238102 473568 238170
rect 473248 238046 473318 238102
rect 473374 238046 473442 238102
rect 473498 238046 473568 238102
rect 473248 237978 473568 238046
rect 473248 237922 473318 237978
rect 473374 237922 473442 237978
rect 473498 237922 473568 237978
rect 473248 237888 473568 237922
rect 503968 238350 504288 238384
rect 503968 238294 504038 238350
rect 504094 238294 504162 238350
rect 504218 238294 504288 238350
rect 503968 238226 504288 238294
rect 503968 238170 504038 238226
rect 504094 238170 504162 238226
rect 504218 238170 504288 238226
rect 503968 238102 504288 238170
rect 503968 238046 504038 238102
rect 504094 238046 504162 238102
rect 504218 238046 504288 238102
rect 503968 237978 504288 238046
rect 503968 237922 504038 237978
rect 504094 237922 504162 237978
rect 504218 237922 504288 237978
rect 503968 237888 504288 237922
rect 534688 238350 535008 238384
rect 534688 238294 534758 238350
rect 534814 238294 534882 238350
rect 534938 238294 535008 238350
rect 534688 238226 535008 238294
rect 534688 238170 534758 238226
rect 534814 238170 534882 238226
rect 534938 238170 535008 238226
rect 534688 238102 535008 238170
rect 534688 238046 534758 238102
rect 534814 238046 534882 238102
rect 534938 238046 535008 238102
rect 534688 237978 535008 238046
rect 534688 237922 534758 237978
rect 534814 237922 534882 237978
rect 534938 237922 535008 237978
rect 534688 237888 535008 237922
rect 565408 238350 565728 238384
rect 565408 238294 565478 238350
rect 565534 238294 565602 238350
rect 565658 238294 565728 238350
rect 565408 238226 565728 238294
rect 565408 238170 565478 238226
rect 565534 238170 565602 238226
rect 565658 238170 565728 238226
rect 565408 238102 565728 238170
rect 565408 238046 565478 238102
rect 565534 238046 565602 238102
rect 565658 238046 565728 238102
rect 565408 237978 565728 238046
rect 565408 237922 565478 237978
rect 565534 237922 565602 237978
rect 565658 237922 565728 237978
rect 565408 237888 565728 237922
rect 585452 232260 585508 271404
rect 585564 253764 585620 284620
rect 589098 274350 589718 291922
rect 589098 274294 589194 274350
rect 589250 274294 589318 274350
rect 589374 274294 589442 274350
rect 589498 274294 589566 274350
rect 589622 274294 589718 274350
rect 589098 274226 589718 274294
rect 589098 274170 589194 274226
rect 589250 274170 589318 274226
rect 589374 274170 589442 274226
rect 589498 274170 589566 274226
rect 589622 274170 589718 274226
rect 589098 274102 589718 274170
rect 589098 274046 589194 274102
rect 589250 274046 589318 274102
rect 589374 274046 589442 274102
rect 589498 274046 589566 274102
rect 589622 274046 589718 274102
rect 589098 273978 589718 274046
rect 589098 273922 589194 273978
rect 589250 273922 589318 273978
rect 589374 273922 589442 273978
rect 589498 273922 589566 273978
rect 589622 273922 589718 273978
rect 585564 253698 585620 253708
rect 587132 258244 587188 258254
rect 585452 232194 585508 232204
rect 6188 228162 6244 228172
rect 585676 231924 585732 231934
rect 27808 226350 28128 226384
rect 27808 226294 27878 226350
rect 27934 226294 28002 226350
rect 28058 226294 28128 226350
rect 27808 226226 28128 226294
rect 27808 226170 27878 226226
rect 27934 226170 28002 226226
rect 28058 226170 28128 226226
rect 27808 226102 28128 226170
rect 27808 226046 27878 226102
rect 27934 226046 28002 226102
rect 28058 226046 28128 226102
rect 27808 225978 28128 226046
rect 27808 225922 27878 225978
rect 27934 225922 28002 225978
rect 28058 225922 28128 225978
rect 27808 225888 28128 225922
rect 58528 226350 58848 226384
rect 58528 226294 58598 226350
rect 58654 226294 58722 226350
rect 58778 226294 58848 226350
rect 58528 226226 58848 226294
rect 58528 226170 58598 226226
rect 58654 226170 58722 226226
rect 58778 226170 58848 226226
rect 58528 226102 58848 226170
rect 58528 226046 58598 226102
rect 58654 226046 58722 226102
rect 58778 226046 58848 226102
rect 58528 225978 58848 226046
rect 58528 225922 58598 225978
rect 58654 225922 58722 225978
rect 58778 225922 58848 225978
rect 58528 225888 58848 225922
rect 89248 226350 89568 226384
rect 89248 226294 89318 226350
rect 89374 226294 89442 226350
rect 89498 226294 89568 226350
rect 89248 226226 89568 226294
rect 89248 226170 89318 226226
rect 89374 226170 89442 226226
rect 89498 226170 89568 226226
rect 89248 226102 89568 226170
rect 89248 226046 89318 226102
rect 89374 226046 89442 226102
rect 89498 226046 89568 226102
rect 89248 225978 89568 226046
rect 89248 225922 89318 225978
rect 89374 225922 89442 225978
rect 89498 225922 89568 225978
rect 89248 225888 89568 225922
rect 119968 226350 120288 226384
rect 119968 226294 120038 226350
rect 120094 226294 120162 226350
rect 120218 226294 120288 226350
rect 119968 226226 120288 226294
rect 119968 226170 120038 226226
rect 120094 226170 120162 226226
rect 120218 226170 120288 226226
rect 119968 226102 120288 226170
rect 119968 226046 120038 226102
rect 120094 226046 120162 226102
rect 120218 226046 120288 226102
rect 119968 225978 120288 226046
rect 119968 225922 120038 225978
rect 120094 225922 120162 225978
rect 120218 225922 120288 225978
rect 119968 225888 120288 225922
rect 150688 226350 151008 226384
rect 150688 226294 150758 226350
rect 150814 226294 150882 226350
rect 150938 226294 151008 226350
rect 150688 226226 151008 226294
rect 150688 226170 150758 226226
rect 150814 226170 150882 226226
rect 150938 226170 151008 226226
rect 150688 226102 151008 226170
rect 150688 226046 150758 226102
rect 150814 226046 150882 226102
rect 150938 226046 151008 226102
rect 150688 225978 151008 226046
rect 150688 225922 150758 225978
rect 150814 225922 150882 225978
rect 150938 225922 151008 225978
rect 150688 225888 151008 225922
rect 181408 226350 181728 226384
rect 181408 226294 181478 226350
rect 181534 226294 181602 226350
rect 181658 226294 181728 226350
rect 181408 226226 181728 226294
rect 181408 226170 181478 226226
rect 181534 226170 181602 226226
rect 181658 226170 181728 226226
rect 181408 226102 181728 226170
rect 181408 226046 181478 226102
rect 181534 226046 181602 226102
rect 181658 226046 181728 226102
rect 181408 225978 181728 226046
rect 181408 225922 181478 225978
rect 181534 225922 181602 225978
rect 181658 225922 181728 225978
rect 181408 225888 181728 225922
rect 212128 226350 212448 226384
rect 212128 226294 212198 226350
rect 212254 226294 212322 226350
rect 212378 226294 212448 226350
rect 212128 226226 212448 226294
rect 212128 226170 212198 226226
rect 212254 226170 212322 226226
rect 212378 226170 212448 226226
rect 212128 226102 212448 226170
rect 212128 226046 212198 226102
rect 212254 226046 212322 226102
rect 212378 226046 212448 226102
rect 212128 225978 212448 226046
rect 212128 225922 212198 225978
rect 212254 225922 212322 225978
rect 212378 225922 212448 225978
rect 212128 225888 212448 225922
rect 242848 226350 243168 226384
rect 242848 226294 242918 226350
rect 242974 226294 243042 226350
rect 243098 226294 243168 226350
rect 242848 226226 243168 226294
rect 242848 226170 242918 226226
rect 242974 226170 243042 226226
rect 243098 226170 243168 226226
rect 242848 226102 243168 226170
rect 242848 226046 242918 226102
rect 242974 226046 243042 226102
rect 243098 226046 243168 226102
rect 242848 225978 243168 226046
rect 242848 225922 242918 225978
rect 242974 225922 243042 225978
rect 243098 225922 243168 225978
rect 242848 225888 243168 225922
rect 273568 226350 273888 226384
rect 273568 226294 273638 226350
rect 273694 226294 273762 226350
rect 273818 226294 273888 226350
rect 273568 226226 273888 226294
rect 273568 226170 273638 226226
rect 273694 226170 273762 226226
rect 273818 226170 273888 226226
rect 273568 226102 273888 226170
rect 273568 226046 273638 226102
rect 273694 226046 273762 226102
rect 273818 226046 273888 226102
rect 273568 225978 273888 226046
rect 273568 225922 273638 225978
rect 273694 225922 273762 225978
rect 273818 225922 273888 225978
rect 273568 225888 273888 225922
rect 304288 226350 304608 226384
rect 304288 226294 304358 226350
rect 304414 226294 304482 226350
rect 304538 226294 304608 226350
rect 304288 226226 304608 226294
rect 304288 226170 304358 226226
rect 304414 226170 304482 226226
rect 304538 226170 304608 226226
rect 304288 226102 304608 226170
rect 304288 226046 304358 226102
rect 304414 226046 304482 226102
rect 304538 226046 304608 226102
rect 304288 225978 304608 226046
rect 304288 225922 304358 225978
rect 304414 225922 304482 225978
rect 304538 225922 304608 225978
rect 304288 225888 304608 225922
rect 335008 226350 335328 226384
rect 335008 226294 335078 226350
rect 335134 226294 335202 226350
rect 335258 226294 335328 226350
rect 335008 226226 335328 226294
rect 335008 226170 335078 226226
rect 335134 226170 335202 226226
rect 335258 226170 335328 226226
rect 335008 226102 335328 226170
rect 335008 226046 335078 226102
rect 335134 226046 335202 226102
rect 335258 226046 335328 226102
rect 335008 225978 335328 226046
rect 335008 225922 335078 225978
rect 335134 225922 335202 225978
rect 335258 225922 335328 225978
rect 335008 225888 335328 225922
rect 365728 226350 366048 226384
rect 365728 226294 365798 226350
rect 365854 226294 365922 226350
rect 365978 226294 366048 226350
rect 365728 226226 366048 226294
rect 365728 226170 365798 226226
rect 365854 226170 365922 226226
rect 365978 226170 366048 226226
rect 365728 226102 366048 226170
rect 365728 226046 365798 226102
rect 365854 226046 365922 226102
rect 365978 226046 366048 226102
rect 365728 225978 366048 226046
rect 365728 225922 365798 225978
rect 365854 225922 365922 225978
rect 365978 225922 366048 225978
rect 365728 225888 366048 225922
rect 396448 226350 396768 226384
rect 396448 226294 396518 226350
rect 396574 226294 396642 226350
rect 396698 226294 396768 226350
rect 396448 226226 396768 226294
rect 396448 226170 396518 226226
rect 396574 226170 396642 226226
rect 396698 226170 396768 226226
rect 396448 226102 396768 226170
rect 396448 226046 396518 226102
rect 396574 226046 396642 226102
rect 396698 226046 396768 226102
rect 396448 225978 396768 226046
rect 396448 225922 396518 225978
rect 396574 225922 396642 225978
rect 396698 225922 396768 225978
rect 396448 225888 396768 225922
rect 427168 226350 427488 226384
rect 427168 226294 427238 226350
rect 427294 226294 427362 226350
rect 427418 226294 427488 226350
rect 427168 226226 427488 226294
rect 427168 226170 427238 226226
rect 427294 226170 427362 226226
rect 427418 226170 427488 226226
rect 427168 226102 427488 226170
rect 427168 226046 427238 226102
rect 427294 226046 427362 226102
rect 427418 226046 427488 226102
rect 427168 225978 427488 226046
rect 427168 225922 427238 225978
rect 427294 225922 427362 225978
rect 427418 225922 427488 225978
rect 427168 225888 427488 225922
rect 457888 226350 458208 226384
rect 457888 226294 457958 226350
rect 458014 226294 458082 226350
rect 458138 226294 458208 226350
rect 457888 226226 458208 226294
rect 457888 226170 457958 226226
rect 458014 226170 458082 226226
rect 458138 226170 458208 226226
rect 457888 226102 458208 226170
rect 457888 226046 457958 226102
rect 458014 226046 458082 226102
rect 458138 226046 458208 226102
rect 457888 225978 458208 226046
rect 457888 225922 457958 225978
rect 458014 225922 458082 225978
rect 458138 225922 458208 225978
rect 457888 225888 458208 225922
rect 488608 226350 488928 226384
rect 488608 226294 488678 226350
rect 488734 226294 488802 226350
rect 488858 226294 488928 226350
rect 488608 226226 488928 226294
rect 488608 226170 488678 226226
rect 488734 226170 488802 226226
rect 488858 226170 488928 226226
rect 488608 226102 488928 226170
rect 488608 226046 488678 226102
rect 488734 226046 488802 226102
rect 488858 226046 488928 226102
rect 488608 225978 488928 226046
rect 488608 225922 488678 225978
rect 488734 225922 488802 225978
rect 488858 225922 488928 225978
rect 488608 225888 488928 225922
rect 519328 226350 519648 226384
rect 519328 226294 519398 226350
rect 519454 226294 519522 226350
rect 519578 226294 519648 226350
rect 519328 226226 519648 226294
rect 519328 226170 519398 226226
rect 519454 226170 519522 226226
rect 519578 226170 519648 226226
rect 519328 226102 519648 226170
rect 519328 226046 519398 226102
rect 519454 226046 519522 226102
rect 519578 226046 519648 226102
rect 519328 225978 519648 226046
rect 519328 225922 519398 225978
rect 519454 225922 519522 225978
rect 519578 225922 519648 225978
rect 519328 225888 519648 225922
rect 550048 226350 550368 226384
rect 550048 226294 550118 226350
rect 550174 226294 550242 226350
rect 550298 226294 550368 226350
rect 550048 226226 550368 226294
rect 550048 226170 550118 226226
rect 550174 226170 550242 226226
rect 550298 226170 550368 226226
rect 550048 226102 550368 226170
rect 550048 226046 550118 226102
rect 550174 226046 550242 226102
rect 550298 226046 550368 226102
rect 550048 225978 550368 226046
rect 550048 225922 550118 225978
rect 550174 225922 550242 225978
rect 550298 225922 550368 225978
rect 550048 225888 550368 225922
rect 5418 220294 5514 220350
rect 5570 220294 5638 220350
rect 5694 220294 5762 220350
rect 5818 220294 5886 220350
rect 5942 220294 6038 220350
rect 5418 220226 6038 220294
rect 12448 220350 12768 220384
rect 12448 220294 12518 220350
rect 12574 220294 12642 220350
rect 12698 220294 12768 220350
rect 5418 220170 5514 220226
rect 5570 220170 5638 220226
rect 5694 220170 5762 220226
rect 5818 220170 5886 220226
rect 5942 220170 6038 220226
rect 5418 220102 6038 220170
rect 5418 220046 5514 220102
rect 5570 220046 5638 220102
rect 5694 220046 5762 220102
rect 5818 220046 5886 220102
rect 5942 220046 6038 220102
rect 5418 219978 6038 220046
rect 5418 219922 5514 219978
rect 5570 219922 5638 219978
rect 5694 219922 5762 219978
rect 5818 219922 5886 219978
rect 5942 219922 6038 219978
rect -956 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 -336 202350
rect -956 202226 -336 202294
rect -956 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 -336 202226
rect -956 202102 -336 202170
rect -956 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 -336 202102
rect -956 201978 -336 202046
rect -956 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 -336 201978
rect -956 184350 -336 201922
rect 5418 202350 6038 219922
rect 6188 220276 6244 220286
rect 6188 207172 6244 220220
rect 12448 220226 12768 220294
rect 12448 220170 12518 220226
rect 12574 220170 12642 220226
rect 12698 220170 12768 220226
rect 12448 220102 12768 220170
rect 12448 220046 12518 220102
rect 12574 220046 12642 220102
rect 12698 220046 12768 220102
rect 12448 219978 12768 220046
rect 12448 219922 12518 219978
rect 12574 219922 12642 219978
rect 12698 219922 12768 219978
rect 12448 219888 12768 219922
rect 43168 220350 43488 220384
rect 43168 220294 43238 220350
rect 43294 220294 43362 220350
rect 43418 220294 43488 220350
rect 43168 220226 43488 220294
rect 43168 220170 43238 220226
rect 43294 220170 43362 220226
rect 43418 220170 43488 220226
rect 43168 220102 43488 220170
rect 43168 220046 43238 220102
rect 43294 220046 43362 220102
rect 43418 220046 43488 220102
rect 43168 219978 43488 220046
rect 43168 219922 43238 219978
rect 43294 219922 43362 219978
rect 43418 219922 43488 219978
rect 43168 219888 43488 219922
rect 73888 220350 74208 220384
rect 73888 220294 73958 220350
rect 74014 220294 74082 220350
rect 74138 220294 74208 220350
rect 73888 220226 74208 220294
rect 73888 220170 73958 220226
rect 74014 220170 74082 220226
rect 74138 220170 74208 220226
rect 73888 220102 74208 220170
rect 73888 220046 73958 220102
rect 74014 220046 74082 220102
rect 74138 220046 74208 220102
rect 73888 219978 74208 220046
rect 73888 219922 73958 219978
rect 74014 219922 74082 219978
rect 74138 219922 74208 219978
rect 73888 219888 74208 219922
rect 104608 220350 104928 220384
rect 104608 220294 104678 220350
rect 104734 220294 104802 220350
rect 104858 220294 104928 220350
rect 104608 220226 104928 220294
rect 104608 220170 104678 220226
rect 104734 220170 104802 220226
rect 104858 220170 104928 220226
rect 104608 220102 104928 220170
rect 104608 220046 104678 220102
rect 104734 220046 104802 220102
rect 104858 220046 104928 220102
rect 104608 219978 104928 220046
rect 104608 219922 104678 219978
rect 104734 219922 104802 219978
rect 104858 219922 104928 219978
rect 104608 219888 104928 219922
rect 135328 220350 135648 220384
rect 135328 220294 135398 220350
rect 135454 220294 135522 220350
rect 135578 220294 135648 220350
rect 135328 220226 135648 220294
rect 135328 220170 135398 220226
rect 135454 220170 135522 220226
rect 135578 220170 135648 220226
rect 135328 220102 135648 220170
rect 135328 220046 135398 220102
rect 135454 220046 135522 220102
rect 135578 220046 135648 220102
rect 135328 219978 135648 220046
rect 135328 219922 135398 219978
rect 135454 219922 135522 219978
rect 135578 219922 135648 219978
rect 135328 219888 135648 219922
rect 166048 220350 166368 220384
rect 166048 220294 166118 220350
rect 166174 220294 166242 220350
rect 166298 220294 166368 220350
rect 166048 220226 166368 220294
rect 166048 220170 166118 220226
rect 166174 220170 166242 220226
rect 166298 220170 166368 220226
rect 166048 220102 166368 220170
rect 166048 220046 166118 220102
rect 166174 220046 166242 220102
rect 166298 220046 166368 220102
rect 166048 219978 166368 220046
rect 166048 219922 166118 219978
rect 166174 219922 166242 219978
rect 166298 219922 166368 219978
rect 166048 219888 166368 219922
rect 196768 220350 197088 220384
rect 196768 220294 196838 220350
rect 196894 220294 196962 220350
rect 197018 220294 197088 220350
rect 196768 220226 197088 220294
rect 196768 220170 196838 220226
rect 196894 220170 196962 220226
rect 197018 220170 197088 220226
rect 196768 220102 197088 220170
rect 196768 220046 196838 220102
rect 196894 220046 196962 220102
rect 197018 220046 197088 220102
rect 196768 219978 197088 220046
rect 196768 219922 196838 219978
rect 196894 219922 196962 219978
rect 197018 219922 197088 219978
rect 196768 219888 197088 219922
rect 227488 220350 227808 220384
rect 227488 220294 227558 220350
rect 227614 220294 227682 220350
rect 227738 220294 227808 220350
rect 227488 220226 227808 220294
rect 227488 220170 227558 220226
rect 227614 220170 227682 220226
rect 227738 220170 227808 220226
rect 227488 220102 227808 220170
rect 227488 220046 227558 220102
rect 227614 220046 227682 220102
rect 227738 220046 227808 220102
rect 227488 219978 227808 220046
rect 227488 219922 227558 219978
rect 227614 219922 227682 219978
rect 227738 219922 227808 219978
rect 227488 219888 227808 219922
rect 258208 220350 258528 220384
rect 258208 220294 258278 220350
rect 258334 220294 258402 220350
rect 258458 220294 258528 220350
rect 258208 220226 258528 220294
rect 258208 220170 258278 220226
rect 258334 220170 258402 220226
rect 258458 220170 258528 220226
rect 258208 220102 258528 220170
rect 258208 220046 258278 220102
rect 258334 220046 258402 220102
rect 258458 220046 258528 220102
rect 258208 219978 258528 220046
rect 258208 219922 258278 219978
rect 258334 219922 258402 219978
rect 258458 219922 258528 219978
rect 258208 219888 258528 219922
rect 288928 220350 289248 220384
rect 288928 220294 288998 220350
rect 289054 220294 289122 220350
rect 289178 220294 289248 220350
rect 288928 220226 289248 220294
rect 288928 220170 288998 220226
rect 289054 220170 289122 220226
rect 289178 220170 289248 220226
rect 288928 220102 289248 220170
rect 288928 220046 288998 220102
rect 289054 220046 289122 220102
rect 289178 220046 289248 220102
rect 288928 219978 289248 220046
rect 288928 219922 288998 219978
rect 289054 219922 289122 219978
rect 289178 219922 289248 219978
rect 288928 219888 289248 219922
rect 319648 220350 319968 220384
rect 319648 220294 319718 220350
rect 319774 220294 319842 220350
rect 319898 220294 319968 220350
rect 319648 220226 319968 220294
rect 319648 220170 319718 220226
rect 319774 220170 319842 220226
rect 319898 220170 319968 220226
rect 319648 220102 319968 220170
rect 319648 220046 319718 220102
rect 319774 220046 319842 220102
rect 319898 220046 319968 220102
rect 319648 219978 319968 220046
rect 319648 219922 319718 219978
rect 319774 219922 319842 219978
rect 319898 219922 319968 219978
rect 319648 219888 319968 219922
rect 350368 220350 350688 220384
rect 350368 220294 350438 220350
rect 350494 220294 350562 220350
rect 350618 220294 350688 220350
rect 350368 220226 350688 220294
rect 350368 220170 350438 220226
rect 350494 220170 350562 220226
rect 350618 220170 350688 220226
rect 350368 220102 350688 220170
rect 350368 220046 350438 220102
rect 350494 220046 350562 220102
rect 350618 220046 350688 220102
rect 350368 219978 350688 220046
rect 350368 219922 350438 219978
rect 350494 219922 350562 219978
rect 350618 219922 350688 219978
rect 350368 219888 350688 219922
rect 381088 220350 381408 220384
rect 381088 220294 381158 220350
rect 381214 220294 381282 220350
rect 381338 220294 381408 220350
rect 381088 220226 381408 220294
rect 381088 220170 381158 220226
rect 381214 220170 381282 220226
rect 381338 220170 381408 220226
rect 381088 220102 381408 220170
rect 381088 220046 381158 220102
rect 381214 220046 381282 220102
rect 381338 220046 381408 220102
rect 381088 219978 381408 220046
rect 381088 219922 381158 219978
rect 381214 219922 381282 219978
rect 381338 219922 381408 219978
rect 381088 219888 381408 219922
rect 411808 220350 412128 220384
rect 411808 220294 411878 220350
rect 411934 220294 412002 220350
rect 412058 220294 412128 220350
rect 411808 220226 412128 220294
rect 411808 220170 411878 220226
rect 411934 220170 412002 220226
rect 412058 220170 412128 220226
rect 411808 220102 412128 220170
rect 411808 220046 411878 220102
rect 411934 220046 412002 220102
rect 412058 220046 412128 220102
rect 411808 219978 412128 220046
rect 411808 219922 411878 219978
rect 411934 219922 412002 219978
rect 412058 219922 412128 219978
rect 411808 219888 412128 219922
rect 442528 220350 442848 220384
rect 442528 220294 442598 220350
rect 442654 220294 442722 220350
rect 442778 220294 442848 220350
rect 442528 220226 442848 220294
rect 442528 220170 442598 220226
rect 442654 220170 442722 220226
rect 442778 220170 442848 220226
rect 442528 220102 442848 220170
rect 442528 220046 442598 220102
rect 442654 220046 442722 220102
rect 442778 220046 442848 220102
rect 442528 219978 442848 220046
rect 442528 219922 442598 219978
rect 442654 219922 442722 219978
rect 442778 219922 442848 219978
rect 442528 219888 442848 219922
rect 473248 220350 473568 220384
rect 473248 220294 473318 220350
rect 473374 220294 473442 220350
rect 473498 220294 473568 220350
rect 473248 220226 473568 220294
rect 473248 220170 473318 220226
rect 473374 220170 473442 220226
rect 473498 220170 473568 220226
rect 473248 220102 473568 220170
rect 473248 220046 473318 220102
rect 473374 220046 473442 220102
rect 473498 220046 473568 220102
rect 473248 219978 473568 220046
rect 473248 219922 473318 219978
rect 473374 219922 473442 219978
rect 473498 219922 473568 219978
rect 473248 219888 473568 219922
rect 503968 220350 504288 220384
rect 503968 220294 504038 220350
rect 504094 220294 504162 220350
rect 504218 220294 504288 220350
rect 503968 220226 504288 220294
rect 503968 220170 504038 220226
rect 504094 220170 504162 220226
rect 504218 220170 504288 220226
rect 503968 220102 504288 220170
rect 503968 220046 504038 220102
rect 504094 220046 504162 220102
rect 504218 220046 504288 220102
rect 503968 219978 504288 220046
rect 503968 219922 504038 219978
rect 504094 219922 504162 219978
rect 504218 219922 504288 219978
rect 503968 219888 504288 219922
rect 534688 220350 535008 220384
rect 534688 220294 534758 220350
rect 534814 220294 534882 220350
rect 534938 220294 535008 220350
rect 534688 220226 535008 220294
rect 534688 220170 534758 220226
rect 534814 220170 534882 220226
rect 534938 220170 535008 220226
rect 534688 220102 535008 220170
rect 534688 220046 534758 220102
rect 534814 220046 534882 220102
rect 534938 220046 535008 220102
rect 534688 219978 535008 220046
rect 534688 219922 534758 219978
rect 534814 219922 534882 219978
rect 534938 219922 535008 219978
rect 534688 219888 535008 219922
rect 565408 220350 565728 220384
rect 565408 220294 565478 220350
rect 565534 220294 565602 220350
rect 565658 220294 565728 220350
rect 565408 220226 565728 220294
rect 565408 220170 565478 220226
rect 565534 220170 565602 220226
rect 565658 220170 565728 220226
rect 565408 220102 565728 220170
rect 565408 220046 565478 220102
rect 565534 220046 565602 220102
rect 565658 220046 565728 220102
rect 565408 219978 565728 220046
rect 565408 219922 565478 219978
rect 565534 219922 565602 219978
rect 565658 219922 565728 219978
rect 565408 219888 565728 219922
rect 585452 218596 585508 218606
rect 27808 208350 28128 208384
rect 27808 208294 27878 208350
rect 27934 208294 28002 208350
rect 28058 208294 28128 208350
rect 27808 208226 28128 208294
rect 27808 208170 27878 208226
rect 27934 208170 28002 208226
rect 28058 208170 28128 208226
rect 27808 208102 28128 208170
rect 27808 208046 27878 208102
rect 27934 208046 28002 208102
rect 28058 208046 28128 208102
rect 27808 207978 28128 208046
rect 27808 207922 27878 207978
rect 27934 207922 28002 207978
rect 28058 207922 28128 207978
rect 27808 207888 28128 207922
rect 58528 208350 58848 208384
rect 58528 208294 58598 208350
rect 58654 208294 58722 208350
rect 58778 208294 58848 208350
rect 58528 208226 58848 208294
rect 58528 208170 58598 208226
rect 58654 208170 58722 208226
rect 58778 208170 58848 208226
rect 58528 208102 58848 208170
rect 58528 208046 58598 208102
rect 58654 208046 58722 208102
rect 58778 208046 58848 208102
rect 58528 207978 58848 208046
rect 58528 207922 58598 207978
rect 58654 207922 58722 207978
rect 58778 207922 58848 207978
rect 58528 207888 58848 207922
rect 89248 208350 89568 208384
rect 89248 208294 89318 208350
rect 89374 208294 89442 208350
rect 89498 208294 89568 208350
rect 89248 208226 89568 208294
rect 89248 208170 89318 208226
rect 89374 208170 89442 208226
rect 89498 208170 89568 208226
rect 89248 208102 89568 208170
rect 89248 208046 89318 208102
rect 89374 208046 89442 208102
rect 89498 208046 89568 208102
rect 89248 207978 89568 208046
rect 89248 207922 89318 207978
rect 89374 207922 89442 207978
rect 89498 207922 89568 207978
rect 89248 207888 89568 207922
rect 119968 208350 120288 208384
rect 119968 208294 120038 208350
rect 120094 208294 120162 208350
rect 120218 208294 120288 208350
rect 119968 208226 120288 208294
rect 119968 208170 120038 208226
rect 120094 208170 120162 208226
rect 120218 208170 120288 208226
rect 119968 208102 120288 208170
rect 119968 208046 120038 208102
rect 120094 208046 120162 208102
rect 120218 208046 120288 208102
rect 119968 207978 120288 208046
rect 119968 207922 120038 207978
rect 120094 207922 120162 207978
rect 120218 207922 120288 207978
rect 119968 207888 120288 207922
rect 150688 208350 151008 208384
rect 150688 208294 150758 208350
rect 150814 208294 150882 208350
rect 150938 208294 151008 208350
rect 150688 208226 151008 208294
rect 150688 208170 150758 208226
rect 150814 208170 150882 208226
rect 150938 208170 151008 208226
rect 150688 208102 151008 208170
rect 150688 208046 150758 208102
rect 150814 208046 150882 208102
rect 150938 208046 151008 208102
rect 150688 207978 151008 208046
rect 150688 207922 150758 207978
rect 150814 207922 150882 207978
rect 150938 207922 151008 207978
rect 150688 207888 151008 207922
rect 181408 208350 181728 208384
rect 181408 208294 181478 208350
rect 181534 208294 181602 208350
rect 181658 208294 181728 208350
rect 181408 208226 181728 208294
rect 181408 208170 181478 208226
rect 181534 208170 181602 208226
rect 181658 208170 181728 208226
rect 181408 208102 181728 208170
rect 181408 208046 181478 208102
rect 181534 208046 181602 208102
rect 181658 208046 181728 208102
rect 181408 207978 181728 208046
rect 181408 207922 181478 207978
rect 181534 207922 181602 207978
rect 181658 207922 181728 207978
rect 181408 207888 181728 207922
rect 212128 208350 212448 208384
rect 212128 208294 212198 208350
rect 212254 208294 212322 208350
rect 212378 208294 212448 208350
rect 212128 208226 212448 208294
rect 212128 208170 212198 208226
rect 212254 208170 212322 208226
rect 212378 208170 212448 208226
rect 212128 208102 212448 208170
rect 212128 208046 212198 208102
rect 212254 208046 212322 208102
rect 212378 208046 212448 208102
rect 212128 207978 212448 208046
rect 212128 207922 212198 207978
rect 212254 207922 212322 207978
rect 212378 207922 212448 207978
rect 212128 207888 212448 207922
rect 242848 208350 243168 208384
rect 242848 208294 242918 208350
rect 242974 208294 243042 208350
rect 243098 208294 243168 208350
rect 242848 208226 243168 208294
rect 242848 208170 242918 208226
rect 242974 208170 243042 208226
rect 243098 208170 243168 208226
rect 242848 208102 243168 208170
rect 242848 208046 242918 208102
rect 242974 208046 243042 208102
rect 243098 208046 243168 208102
rect 242848 207978 243168 208046
rect 242848 207922 242918 207978
rect 242974 207922 243042 207978
rect 243098 207922 243168 207978
rect 242848 207888 243168 207922
rect 273568 208350 273888 208384
rect 273568 208294 273638 208350
rect 273694 208294 273762 208350
rect 273818 208294 273888 208350
rect 273568 208226 273888 208294
rect 273568 208170 273638 208226
rect 273694 208170 273762 208226
rect 273818 208170 273888 208226
rect 273568 208102 273888 208170
rect 273568 208046 273638 208102
rect 273694 208046 273762 208102
rect 273818 208046 273888 208102
rect 273568 207978 273888 208046
rect 273568 207922 273638 207978
rect 273694 207922 273762 207978
rect 273818 207922 273888 207978
rect 273568 207888 273888 207922
rect 304288 208350 304608 208384
rect 304288 208294 304358 208350
rect 304414 208294 304482 208350
rect 304538 208294 304608 208350
rect 304288 208226 304608 208294
rect 304288 208170 304358 208226
rect 304414 208170 304482 208226
rect 304538 208170 304608 208226
rect 304288 208102 304608 208170
rect 304288 208046 304358 208102
rect 304414 208046 304482 208102
rect 304538 208046 304608 208102
rect 304288 207978 304608 208046
rect 304288 207922 304358 207978
rect 304414 207922 304482 207978
rect 304538 207922 304608 207978
rect 304288 207888 304608 207922
rect 335008 208350 335328 208384
rect 335008 208294 335078 208350
rect 335134 208294 335202 208350
rect 335258 208294 335328 208350
rect 335008 208226 335328 208294
rect 335008 208170 335078 208226
rect 335134 208170 335202 208226
rect 335258 208170 335328 208226
rect 335008 208102 335328 208170
rect 335008 208046 335078 208102
rect 335134 208046 335202 208102
rect 335258 208046 335328 208102
rect 335008 207978 335328 208046
rect 335008 207922 335078 207978
rect 335134 207922 335202 207978
rect 335258 207922 335328 207978
rect 335008 207888 335328 207922
rect 365728 208350 366048 208384
rect 365728 208294 365798 208350
rect 365854 208294 365922 208350
rect 365978 208294 366048 208350
rect 365728 208226 366048 208294
rect 365728 208170 365798 208226
rect 365854 208170 365922 208226
rect 365978 208170 366048 208226
rect 365728 208102 366048 208170
rect 365728 208046 365798 208102
rect 365854 208046 365922 208102
rect 365978 208046 366048 208102
rect 365728 207978 366048 208046
rect 365728 207922 365798 207978
rect 365854 207922 365922 207978
rect 365978 207922 366048 207978
rect 365728 207888 366048 207922
rect 396448 208350 396768 208384
rect 396448 208294 396518 208350
rect 396574 208294 396642 208350
rect 396698 208294 396768 208350
rect 396448 208226 396768 208294
rect 396448 208170 396518 208226
rect 396574 208170 396642 208226
rect 396698 208170 396768 208226
rect 396448 208102 396768 208170
rect 396448 208046 396518 208102
rect 396574 208046 396642 208102
rect 396698 208046 396768 208102
rect 396448 207978 396768 208046
rect 396448 207922 396518 207978
rect 396574 207922 396642 207978
rect 396698 207922 396768 207978
rect 396448 207888 396768 207922
rect 427168 208350 427488 208384
rect 427168 208294 427238 208350
rect 427294 208294 427362 208350
rect 427418 208294 427488 208350
rect 427168 208226 427488 208294
rect 427168 208170 427238 208226
rect 427294 208170 427362 208226
rect 427418 208170 427488 208226
rect 427168 208102 427488 208170
rect 427168 208046 427238 208102
rect 427294 208046 427362 208102
rect 427418 208046 427488 208102
rect 427168 207978 427488 208046
rect 427168 207922 427238 207978
rect 427294 207922 427362 207978
rect 427418 207922 427488 207978
rect 427168 207888 427488 207922
rect 457888 208350 458208 208384
rect 457888 208294 457958 208350
rect 458014 208294 458082 208350
rect 458138 208294 458208 208350
rect 457888 208226 458208 208294
rect 457888 208170 457958 208226
rect 458014 208170 458082 208226
rect 458138 208170 458208 208226
rect 457888 208102 458208 208170
rect 457888 208046 457958 208102
rect 458014 208046 458082 208102
rect 458138 208046 458208 208102
rect 457888 207978 458208 208046
rect 457888 207922 457958 207978
rect 458014 207922 458082 207978
rect 458138 207922 458208 207978
rect 457888 207888 458208 207922
rect 488608 208350 488928 208384
rect 488608 208294 488678 208350
rect 488734 208294 488802 208350
rect 488858 208294 488928 208350
rect 488608 208226 488928 208294
rect 488608 208170 488678 208226
rect 488734 208170 488802 208226
rect 488858 208170 488928 208226
rect 488608 208102 488928 208170
rect 488608 208046 488678 208102
rect 488734 208046 488802 208102
rect 488858 208046 488928 208102
rect 488608 207978 488928 208046
rect 488608 207922 488678 207978
rect 488734 207922 488802 207978
rect 488858 207922 488928 207978
rect 488608 207888 488928 207922
rect 519328 208350 519648 208384
rect 519328 208294 519398 208350
rect 519454 208294 519522 208350
rect 519578 208294 519648 208350
rect 519328 208226 519648 208294
rect 519328 208170 519398 208226
rect 519454 208170 519522 208226
rect 519578 208170 519648 208226
rect 519328 208102 519648 208170
rect 519328 208046 519398 208102
rect 519454 208046 519522 208102
rect 519578 208046 519648 208102
rect 519328 207978 519648 208046
rect 519328 207922 519398 207978
rect 519454 207922 519522 207978
rect 519578 207922 519648 207978
rect 519328 207888 519648 207922
rect 550048 208350 550368 208384
rect 550048 208294 550118 208350
rect 550174 208294 550242 208350
rect 550298 208294 550368 208350
rect 550048 208226 550368 208294
rect 550048 208170 550118 208226
rect 550174 208170 550242 208226
rect 550298 208170 550368 208226
rect 550048 208102 550368 208170
rect 550048 208046 550118 208102
rect 550174 208046 550242 208102
rect 550298 208046 550368 208102
rect 550048 207978 550368 208046
rect 550048 207922 550118 207978
rect 550174 207922 550242 207978
rect 550298 207922 550368 207978
rect 550048 207888 550368 207922
rect 6188 207106 6244 207116
rect 5418 202294 5514 202350
rect 5570 202294 5638 202350
rect 5694 202294 5762 202350
rect 5818 202294 5886 202350
rect 5942 202294 6038 202350
rect 5418 202226 6038 202294
rect 5418 202170 5514 202226
rect 5570 202170 5638 202226
rect 5694 202170 5762 202226
rect 5818 202170 5886 202226
rect 5942 202170 6038 202226
rect 5418 202102 6038 202170
rect 5418 202046 5514 202102
rect 5570 202046 5638 202102
rect 5694 202046 5762 202102
rect 5818 202046 5886 202102
rect 5942 202046 6038 202102
rect 5418 201978 6038 202046
rect 5418 201922 5514 201978
rect 5570 201922 5638 201978
rect 5694 201922 5762 201978
rect 5818 201922 5886 201978
rect 5942 201922 6038 201978
rect -956 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 -336 184350
rect -956 184226 -336 184294
rect -956 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 -336 184226
rect -956 184102 -336 184170
rect -956 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 -336 184102
rect -956 183978 -336 184046
rect -956 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 -336 183978
rect -956 166350 -336 183922
rect 4172 192052 4228 192062
rect 4172 175588 4228 191996
rect 5418 184350 6038 201922
rect 6188 206164 6244 206174
rect 6188 186116 6244 206108
rect 12448 202350 12768 202384
rect 12448 202294 12518 202350
rect 12574 202294 12642 202350
rect 12698 202294 12768 202350
rect 12448 202226 12768 202294
rect 12448 202170 12518 202226
rect 12574 202170 12642 202226
rect 12698 202170 12768 202226
rect 12448 202102 12768 202170
rect 12448 202046 12518 202102
rect 12574 202046 12642 202102
rect 12698 202046 12768 202102
rect 12448 201978 12768 202046
rect 12448 201922 12518 201978
rect 12574 201922 12642 201978
rect 12698 201922 12768 201978
rect 12448 201888 12768 201922
rect 43168 202350 43488 202384
rect 43168 202294 43238 202350
rect 43294 202294 43362 202350
rect 43418 202294 43488 202350
rect 43168 202226 43488 202294
rect 43168 202170 43238 202226
rect 43294 202170 43362 202226
rect 43418 202170 43488 202226
rect 43168 202102 43488 202170
rect 43168 202046 43238 202102
rect 43294 202046 43362 202102
rect 43418 202046 43488 202102
rect 43168 201978 43488 202046
rect 43168 201922 43238 201978
rect 43294 201922 43362 201978
rect 43418 201922 43488 201978
rect 43168 201888 43488 201922
rect 73888 202350 74208 202384
rect 73888 202294 73958 202350
rect 74014 202294 74082 202350
rect 74138 202294 74208 202350
rect 73888 202226 74208 202294
rect 73888 202170 73958 202226
rect 74014 202170 74082 202226
rect 74138 202170 74208 202226
rect 73888 202102 74208 202170
rect 73888 202046 73958 202102
rect 74014 202046 74082 202102
rect 74138 202046 74208 202102
rect 73888 201978 74208 202046
rect 73888 201922 73958 201978
rect 74014 201922 74082 201978
rect 74138 201922 74208 201978
rect 73888 201888 74208 201922
rect 104608 202350 104928 202384
rect 104608 202294 104678 202350
rect 104734 202294 104802 202350
rect 104858 202294 104928 202350
rect 104608 202226 104928 202294
rect 104608 202170 104678 202226
rect 104734 202170 104802 202226
rect 104858 202170 104928 202226
rect 104608 202102 104928 202170
rect 104608 202046 104678 202102
rect 104734 202046 104802 202102
rect 104858 202046 104928 202102
rect 104608 201978 104928 202046
rect 104608 201922 104678 201978
rect 104734 201922 104802 201978
rect 104858 201922 104928 201978
rect 104608 201888 104928 201922
rect 135328 202350 135648 202384
rect 135328 202294 135398 202350
rect 135454 202294 135522 202350
rect 135578 202294 135648 202350
rect 135328 202226 135648 202294
rect 135328 202170 135398 202226
rect 135454 202170 135522 202226
rect 135578 202170 135648 202226
rect 135328 202102 135648 202170
rect 135328 202046 135398 202102
rect 135454 202046 135522 202102
rect 135578 202046 135648 202102
rect 135328 201978 135648 202046
rect 135328 201922 135398 201978
rect 135454 201922 135522 201978
rect 135578 201922 135648 201978
rect 135328 201888 135648 201922
rect 166048 202350 166368 202384
rect 166048 202294 166118 202350
rect 166174 202294 166242 202350
rect 166298 202294 166368 202350
rect 166048 202226 166368 202294
rect 166048 202170 166118 202226
rect 166174 202170 166242 202226
rect 166298 202170 166368 202226
rect 166048 202102 166368 202170
rect 166048 202046 166118 202102
rect 166174 202046 166242 202102
rect 166298 202046 166368 202102
rect 166048 201978 166368 202046
rect 166048 201922 166118 201978
rect 166174 201922 166242 201978
rect 166298 201922 166368 201978
rect 166048 201888 166368 201922
rect 196768 202350 197088 202384
rect 196768 202294 196838 202350
rect 196894 202294 196962 202350
rect 197018 202294 197088 202350
rect 196768 202226 197088 202294
rect 196768 202170 196838 202226
rect 196894 202170 196962 202226
rect 197018 202170 197088 202226
rect 196768 202102 197088 202170
rect 196768 202046 196838 202102
rect 196894 202046 196962 202102
rect 197018 202046 197088 202102
rect 196768 201978 197088 202046
rect 196768 201922 196838 201978
rect 196894 201922 196962 201978
rect 197018 201922 197088 201978
rect 196768 201888 197088 201922
rect 227488 202350 227808 202384
rect 227488 202294 227558 202350
rect 227614 202294 227682 202350
rect 227738 202294 227808 202350
rect 227488 202226 227808 202294
rect 227488 202170 227558 202226
rect 227614 202170 227682 202226
rect 227738 202170 227808 202226
rect 227488 202102 227808 202170
rect 227488 202046 227558 202102
rect 227614 202046 227682 202102
rect 227738 202046 227808 202102
rect 227488 201978 227808 202046
rect 227488 201922 227558 201978
rect 227614 201922 227682 201978
rect 227738 201922 227808 201978
rect 227488 201888 227808 201922
rect 258208 202350 258528 202384
rect 258208 202294 258278 202350
rect 258334 202294 258402 202350
rect 258458 202294 258528 202350
rect 258208 202226 258528 202294
rect 258208 202170 258278 202226
rect 258334 202170 258402 202226
rect 258458 202170 258528 202226
rect 258208 202102 258528 202170
rect 258208 202046 258278 202102
rect 258334 202046 258402 202102
rect 258458 202046 258528 202102
rect 258208 201978 258528 202046
rect 258208 201922 258278 201978
rect 258334 201922 258402 201978
rect 258458 201922 258528 201978
rect 258208 201888 258528 201922
rect 288928 202350 289248 202384
rect 288928 202294 288998 202350
rect 289054 202294 289122 202350
rect 289178 202294 289248 202350
rect 288928 202226 289248 202294
rect 288928 202170 288998 202226
rect 289054 202170 289122 202226
rect 289178 202170 289248 202226
rect 288928 202102 289248 202170
rect 288928 202046 288998 202102
rect 289054 202046 289122 202102
rect 289178 202046 289248 202102
rect 288928 201978 289248 202046
rect 288928 201922 288998 201978
rect 289054 201922 289122 201978
rect 289178 201922 289248 201978
rect 288928 201888 289248 201922
rect 319648 202350 319968 202384
rect 319648 202294 319718 202350
rect 319774 202294 319842 202350
rect 319898 202294 319968 202350
rect 319648 202226 319968 202294
rect 319648 202170 319718 202226
rect 319774 202170 319842 202226
rect 319898 202170 319968 202226
rect 319648 202102 319968 202170
rect 319648 202046 319718 202102
rect 319774 202046 319842 202102
rect 319898 202046 319968 202102
rect 319648 201978 319968 202046
rect 319648 201922 319718 201978
rect 319774 201922 319842 201978
rect 319898 201922 319968 201978
rect 319648 201888 319968 201922
rect 350368 202350 350688 202384
rect 350368 202294 350438 202350
rect 350494 202294 350562 202350
rect 350618 202294 350688 202350
rect 350368 202226 350688 202294
rect 350368 202170 350438 202226
rect 350494 202170 350562 202226
rect 350618 202170 350688 202226
rect 350368 202102 350688 202170
rect 350368 202046 350438 202102
rect 350494 202046 350562 202102
rect 350618 202046 350688 202102
rect 350368 201978 350688 202046
rect 350368 201922 350438 201978
rect 350494 201922 350562 201978
rect 350618 201922 350688 201978
rect 350368 201888 350688 201922
rect 381088 202350 381408 202384
rect 381088 202294 381158 202350
rect 381214 202294 381282 202350
rect 381338 202294 381408 202350
rect 381088 202226 381408 202294
rect 381088 202170 381158 202226
rect 381214 202170 381282 202226
rect 381338 202170 381408 202226
rect 381088 202102 381408 202170
rect 381088 202046 381158 202102
rect 381214 202046 381282 202102
rect 381338 202046 381408 202102
rect 381088 201978 381408 202046
rect 381088 201922 381158 201978
rect 381214 201922 381282 201978
rect 381338 201922 381408 201978
rect 381088 201888 381408 201922
rect 411808 202350 412128 202384
rect 411808 202294 411878 202350
rect 411934 202294 412002 202350
rect 412058 202294 412128 202350
rect 411808 202226 412128 202294
rect 411808 202170 411878 202226
rect 411934 202170 412002 202226
rect 412058 202170 412128 202226
rect 411808 202102 412128 202170
rect 411808 202046 411878 202102
rect 411934 202046 412002 202102
rect 412058 202046 412128 202102
rect 411808 201978 412128 202046
rect 411808 201922 411878 201978
rect 411934 201922 412002 201978
rect 412058 201922 412128 201978
rect 411808 201888 412128 201922
rect 442528 202350 442848 202384
rect 442528 202294 442598 202350
rect 442654 202294 442722 202350
rect 442778 202294 442848 202350
rect 442528 202226 442848 202294
rect 442528 202170 442598 202226
rect 442654 202170 442722 202226
rect 442778 202170 442848 202226
rect 442528 202102 442848 202170
rect 442528 202046 442598 202102
rect 442654 202046 442722 202102
rect 442778 202046 442848 202102
rect 442528 201978 442848 202046
rect 442528 201922 442598 201978
rect 442654 201922 442722 201978
rect 442778 201922 442848 201978
rect 442528 201888 442848 201922
rect 473248 202350 473568 202384
rect 473248 202294 473318 202350
rect 473374 202294 473442 202350
rect 473498 202294 473568 202350
rect 473248 202226 473568 202294
rect 473248 202170 473318 202226
rect 473374 202170 473442 202226
rect 473498 202170 473568 202226
rect 473248 202102 473568 202170
rect 473248 202046 473318 202102
rect 473374 202046 473442 202102
rect 473498 202046 473568 202102
rect 473248 201978 473568 202046
rect 473248 201922 473318 201978
rect 473374 201922 473442 201978
rect 473498 201922 473568 201978
rect 473248 201888 473568 201922
rect 503968 202350 504288 202384
rect 503968 202294 504038 202350
rect 504094 202294 504162 202350
rect 504218 202294 504288 202350
rect 503968 202226 504288 202294
rect 503968 202170 504038 202226
rect 504094 202170 504162 202226
rect 504218 202170 504288 202226
rect 503968 202102 504288 202170
rect 503968 202046 504038 202102
rect 504094 202046 504162 202102
rect 504218 202046 504288 202102
rect 503968 201978 504288 202046
rect 503968 201922 504038 201978
rect 504094 201922 504162 201978
rect 504218 201922 504288 201978
rect 503968 201888 504288 201922
rect 534688 202350 535008 202384
rect 534688 202294 534758 202350
rect 534814 202294 534882 202350
rect 534938 202294 535008 202350
rect 534688 202226 535008 202294
rect 534688 202170 534758 202226
rect 534814 202170 534882 202226
rect 534938 202170 535008 202226
rect 534688 202102 535008 202170
rect 534688 202046 534758 202102
rect 534814 202046 534882 202102
rect 534938 202046 535008 202102
rect 534688 201978 535008 202046
rect 534688 201922 534758 201978
rect 534814 201922 534882 201978
rect 534938 201922 535008 201978
rect 534688 201888 535008 201922
rect 565408 202350 565728 202384
rect 565408 202294 565478 202350
rect 565534 202294 565602 202350
rect 565658 202294 565728 202350
rect 565408 202226 565728 202294
rect 565408 202170 565478 202226
rect 565534 202170 565602 202226
rect 565658 202170 565728 202226
rect 565408 202102 565728 202170
rect 565408 202046 565478 202102
rect 565534 202046 565602 202102
rect 565658 202046 565728 202102
rect 565408 201978 565728 202046
rect 565408 201922 565478 201978
rect 565534 201922 565602 201978
rect 565658 201922 565728 201978
rect 565408 201888 565728 201922
rect 27808 190350 28128 190384
rect 27808 190294 27878 190350
rect 27934 190294 28002 190350
rect 28058 190294 28128 190350
rect 27808 190226 28128 190294
rect 27808 190170 27878 190226
rect 27934 190170 28002 190226
rect 28058 190170 28128 190226
rect 27808 190102 28128 190170
rect 27808 190046 27878 190102
rect 27934 190046 28002 190102
rect 28058 190046 28128 190102
rect 27808 189978 28128 190046
rect 27808 189922 27878 189978
rect 27934 189922 28002 189978
rect 28058 189922 28128 189978
rect 27808 189888 28128 189922
rect 58528 190350 58848 190384
rect 58528 190294 58598 190350
rect 58654 190294 58722 190350
rect 58778 190294 58848 190350
rect 58528 190226 58848 190294
rect 58528 190170 58598 190226
rect 58654 190170 58722 190226
rect 58778 190170 58848 190226
rect 58528 190102 58848 190170
rect 58528 190046 58598 190102
rect 58654 190046 58722 190102
rect 58778 190046 58848 190102
rect 58528 189978 58848 190046
rect 58528 189922 58598 189978
rect 58654 189922 58722 189978
rect 58778 189922 58848 189978
rect 58528 189888 58848 189922
rect 89248 190350 89568 190384
rect 89248 190294 89318 190350
rect 89374 190294 89442 190350
rect 89498 190294 89568 190350
rect 89248 190226 89568 190294
rect 89248 190170 89318 190226
rect 89374 190170 89442 190226
rect 89498 190170 89568 190226
rect 89248 190102 89568 190170
rect 89248 190046 89318 190102
rect 89374 190046 89442 190102
rect 89498 190046 89568 190102
rect 89248 189978 89568 190046
rect 89248 189922 89318 189978
rect 89374 189922 89442 189978
rect 89498 189922 89568 189978
rect 89248 189888 89568 189922
rect 119968 190350 120288 190384
rect 119968 190294 120038 190350
rect 120094 190294 120162 190350
rect 120218 190294 120288 190350
rect 119968 190226 120288 190294
rect 119968 190170 120038 190226
rect 120094 190170 120162 190226
rect 120218 190170 120288 190226
rect 119968 190102 120288 190170
rect 119968 190046 120038 190102
rect 120094 190046 120162 190102
rect 120218 190046 120288 190102
rect 119968 189978 120288 190046
rect 119968 189922 120038 189978
rect 120094 189922 120162 189978
rect 120218 189922 120288 189978
rect 119968 189888 120288 189922
rect 150688 190350 151008 190384
rect 150688 190294 150758 190350
rect 150814 190294 150882 190350
rect 150938 190294 151008 190350
rect 150688 190226 151008 190294
rect 150688 190170 150758 190226
rect 150814 190170 150882 190226
rect 150938 190170 151008 190226
rect 150688 190102 151008 190170
rect 150688 190046 150758 190102
rect 150814 190046 150882 190102
rect 150938 190046 151008 190102
rect 150688 189978 151008 190046
rect 150688 189922 150758 189978
rect 150814 189922 150882 189978
rect 150938 189922 151008 189978
rect 150688 189888 151008 189922
rect 181408 190350 181728 190384
rect 181408 190294 181478 190350
rect 181534 190294 181602 190350
rect 181658 190294 181728 190350
rect 181408 190226 181728 190294
rect 181408 190170 181478 190226
rect 181534 190170 181602 190226
rect 181658 190170 181728 190226
rect 181408 190102 181728 190170
rect 181408 190046 181478 190102
rect 181534 190046 181602 190102
rect 181658 190046 181728 190102
rect 181408 189978 181728 190046
rect 181408 189922 181478 189978
rect 181534 189922 181602 189978
rect 181658 189922 181728 189978
rect 181408 189888 181728 189922
rect 212128 190350 212448 190384
rect 212128 190294 212198 190350
rect 212254 190294 212322 190350
rect 212378 190294 212448 190350
rect 212128 190226 212448 190294
rect 212128 190170 212198 190226
rect 212254 190170 212322 190226
rect 212378 190170 212448 190226
rect 212128 190102 212448 190170
rect 212128 190046 212198 190102
rect 212254 190046 212322 190102
rect 212378 190046 212448 190102
rect 212128 189978 212448 190046
rect 212128 189922 212198 189978
rect 212254 189922 212322 189978
rect 212378 189922 212448 189978
rect 212128 189888 212448 189922
rect 242848 190350 243168 190384
rect 242848 190294 242918 190350
rect 242974 190294 243042 190350
rect 243098 190294 243168 190350
rect 242848 190226 243168 190294
rect 242848 190170 242918 190226
rect 242974 190170 243042 190226
rect 243098 190170 243168 190226
rect 242848 190102 243168 190170
rect 242848 190046 242918 190102
rect 242974 190046 243042 190102
rect 243098 190046 243168 190102
rect 242848 189978 243168 190046
rect 242848 189922 242918 189978
rect 242974 189922 243042 189978
rect 243098 189922 243168 189978
rect 242848 189888 243168 189922
rect 273568 190350 273888 190384
rect 273568 190294 273638 190350
rect 273694 190294 273762 190350
rect 273818 190294 273888 190350
rect 273568 190226 273888 190294
rect 273568 190170 273638 190226
rect 273694 190170 273762 190226
rect 273818 190170 273888 190226
rect 273568 190102 273888 190170
rect 273568 190046 273638 190102
rect 273694 190046 273762 190102
rect 273818 190046 273888 190102
rect 273568 189978 273888 190046
rect 273568 189922 273638 189978
rect 273694 189922 273762 189978
rect 273818 189922 273888 189978
rect 273568 189888 273888 189922
rect 304288 190350 304608 190384
rect 304288 190294 304358 190350
rect 304414 190294 304482 190350
rect 304538 190294 304608 190350
rect 304288 190226 304608 190294
rect 304288 190170 304358 190226
rect 304414 190170 304482 190226
rect 304538 190170 304608 190226
rect 304288 190102 304608 190170
rect 304288 190046 304358 190102
rect 304414 190046 304482 190102
rect 304538 190046 304608 190102
rect 304288 189978 304608 190046
rect 304288 189922 304358 189978
rect 304414 189922 304482 189978
rect 304538 189922 304608 189978
rect 304288 189888 304608 189922
rect 335008 190350 335328 190384
rect 335008 190294 335078 190350
rect 335134 190294 335202 190350
rect 335258 190294 335328 190350
rect 335008 190226 335328 190294
rect 335008 190170 335078 190226
rect 335134 190170 335202 190226
rect 335258 190170 335328 190226
rect 335008 190102 335328 190170
rect 335008 190046 335078 190102
rect 335134 190046 335202 190102
rect 335258 190046 335328 190102
rect 335008 189978 335328 190046
rect 335008 189922 335078 189978
rect 335134 189922 335202 189978
rect 335258 189922 335328 189978
rect 335008 189888 335328 189922
rect 365728 190350 366048 190384
rect 365728 190294 365798 190350
rect 365854 190294 365922 190350
rect 365978 190294 366048 190350
rect 365728 190226 366048 190294
rect 365728 190170 365798 190226
rect 365854 190170 365922 190226
rect 365978 190170 366048 190226
rect 365728 190102 366048 190170
rect 365728 190046 365798 190102
rect 365854 190046 365922 190102
rect 365978 190046 366048 190102
rect 365728 189978 366048 190046
rect 365728 189922 365798 189978
rect 365854 189922 365922 189978
rect 365978 189922 366048 189978
rect 365728 189888 366048 189922
rect 396448 190350 396768 190384
rect 396448 190294 396518 190350
rect 396574 190294 396642 190350
rect 396698 190294 396768 190350
rect 396448 190226 396768 190294
rect 396448 190170 396518 190226
rect 396574 190170 396642 190226
rect 396698 190170 396768 190226
rect 396448 190102 396768 190170
rect 396448 190046 396518 190102
rect 396574 190046 396642 190102
rect 396698 190046 396768 190102
rect 396448 189978 396768 190046
rect 396448 189922 396518 189978
rect 396574 189922 396642 189978
rect 396698 189922 396768 189978
rect 396448 189888 396768 189922
rect 427168 190350 427488 190384
rect 427168 190294 427238 190350
rect 427294 190294 427362 190350
rect 427418 190294 427488 190350
rect 427168 190226 427488 190294
rect 427168 190170 427238 190226
rect 427294 190170 427362 190226
rect 427418 190170 427488 190226
rect 427168 190102 427488 190170
rect 427168 190046 427238 190102
rect 427294 190046 427362 190102
rect 427418 190046 427488 190102
rect 427168 189978 427488 190046
rect 427168 189922 427238 189978
rect 427294 189922 427362 189978
rect 427418 189922 427488 189978
rect 427168 189888 427488 189922
rect 457888 190350 458208 190384
rect 457888 190294 457958 190350
rect 458014 190294 458082 190350
rect 458138 190294 458208 190350
rect 457888 190226 458208 190294
rect 457888 190170 457958 190226
rect 458014 190170 458082 190226
rect 458138 190170 458208 190226
rect 457888 190102 458208 190170
rect 457888 190046 457958 190102
rect 458014 190046 458082 190102
rect 458138 190046 458208 190102
rect 457888 189978 458208 190046
rect 457888 189922 457958 189978
rect 458014 189922 458082 189978
rect 458138 189922 458208 189978
rect 457888 189888 458208 189922
rect 488608 190350 488928 190384
rect 488608 190294 488678 190350
rect 488734 190294 488802 190350
rect 488858 190294 488928 190350
rect 488608 190226 488928 190294
rect 488608 190170 488678 190226
rect 488734 190170 488802 190226
rect 488858 190170 488928 190226
rect 488608 190102 488928 190170
rect 488608 190046 488678 190102
rect 488734 190046 488802 190102
rect 488858 190046 488928 190102
rect 488608 189978 488928 190046
rect 488608 189922 488678 189978
rect 488734 189922 488802 189978
rect 488858 189922 488928 189978
rect 488608 189888 488928 189922
rect 519328 190350 519648 190384
rect 519328 190294 519398 190350
rect 519454 190294 519522 190350
rect 519578 190294 519648 190350
rect 519328 190226 519648 190294
rect 519328 190170 519398 190226
rect 519454 190170 519522 190226
rect 519578 190170 519648 190226
rect 519328 190102 519648 190170
rect 519328 190046 519398 190102
rect 519454 190046 519522 190102
rect 519578 190046 519648 190102
rect 519328 189978 519648 190046
rect 519328 189922 519398 189978
rect 519454 189922 519522 189978
rect 519578 189922 519648 189978
rect 519328 189888 519648 189922
rect 550048 190350 550368 190384
rect 550048 190294 550118 190350
rect 550174 190294 550242 190350
rect 550298 190294 550368 190350
rect 550048 190226 550368 190294
rect 550048 190170 550118 190226
rect 550174 190170 550242 190226
rect 550298 190170 550368 190226
rect 550048 190102 550368 190170
rect 550048 190046 550118 190102
rect 550174 190046 550242 190102
rect 550298 190046 550368 190102
rect 550048 189978 550368 190046
rect 550048 189922 550118 189978
rect 550174 189922 550242 189978
rect 550298 189922 550368 189978
rect 550048 189888 550368 189922
rect 585452 189252 585508 218540
rect 585452 189186 585508 189196
rect 585564 205380 585620 205390
rect 6188 186050 6244 186060
rect 5418 184294 5514 184350
rect 5570 184294 5638 184350
rect 5694 184294 5762 184350
rect 5818 184294 5886 184350
rect 5942 184294 6038 184350
rect 5418 184226 6038 184294
rect 5418 184170 5514 184226
rect 5570 184170 5638 184226
rect 5694 184170 5762 184226
rect 5818 184170 5886 184226
rect 5942 184170 6038 184226
rect 5418 184102 6038 184170
rect 5418 184046 5514 184102
rect 5570 184046 5638 184102
rect 5694 184046 5762 184102
rect 5818 184046 5886 184102
rect 5942 184046 6038 184102
rect 5418 183978 6038 184046
rect 5418 183922 5514 183978
rect 5570 183922 5638 183978
rect 5694 183922 5762 183978
rect 5818 183922 5886 183978
rect 5942 183922 6038 183978
rect 4172 175522 4228 175532
rect 4284 177940 4340 177950
rect -956 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 -336 166350
rect -956 166226 -336 166294
rect -956 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 -336 166226
rect -956 166102 -336 166170
rect -956 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 -336 166102
rect -956 165978 -336 166046
rect -956 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 -336 165978
rect -956 148350 -336 165922
rect 4284 165060 4340 177884
rect 4284 164994 4340 165004
rect 5418 166350 6038 183922
rect 12448 184350 12768 184384
rect 12448 184294 12518 184350
rect 12574 184294 12642 184350
rect 12698 184294 12768 184350
rect 12448 184226 12768 184294
rect 12448 184170 12518 184226
rect 12574 184170 12642 184226
rect 12698 184170 12768 184226
rect 12448 184102 12768 184170
rect 12448 184046 12518 184102
rect 12574 184046 12642 184102
rect 12698 184046 12768 184102
rect 12448 183978 12768 184046
rect 12448 183922 12518 183978
rect 12574 183922 12642 183978
rect 12698 183922 12768 183978
rect 12448 183888 12768 183922
rect 43168 184350 43488 184384
rect 43168 184294 43238 184350
rect 43294 184294 43362 184350
rect 43418 184294 43488 184350
rect 43168 184226 43488 184294
rect 43168 184170 43238 184226
rect 43294 184170 43362 184226
rect 43418 184170 43488 184226
rect 43168 184102 43488 184170
rect 43168 184046 43238 184102
rect 43294 184046 43362 184102
rect 43418 184046 43488 184102
rect 43168 183978 43488 184046
rect 43168 183922 43238 183978
rect 43294 183922 43362 183978
rect 43418 183922 43488 183978
rect 43168 183888 43488 183922
rect 73888 184350 74208 184384
rect 73888 184294 73958 184350
rect 74014 184294 74082 184350
rect 74138 184294 74208 184350
rect 73888 184226 74208 184294
rect 73888 184170 73958 184226
rect 74014 184170 74082 184226
rect 74138 184170 74208 184226
rect 73888 184102 74208 184170
rect 73888 184046 73958 184102
rect 74014 184046 74082 184102
rect 74138 184046 74208 184102
rect 73888 183978 74208 184046
rect 73888 183922 73958 183978
rect 74014 183922 74082 183978
rect 74138 183922 74208 183978
rect 73888 183888 74208 183922
rect 104608 184350 104928 184384
rect 104608 184294 104678 184350
rect 104734 184294 104802 184350
rect 104858 184294 104928 184350
rect 104608 184226 104928 184294
rect 104608 184170 104678 184226
rect 104734 184170 104802 184226
rect 104858 184170 104928 184226
rect 104608 184102 104928 184170
rect 104608 184046 104678 184102
rect 104734 184046 104802 184102
rect 104858 184046 104928 184102
rect 104608 183978 104928 184046
rect 104608 183922 104678 183978
rect 104734 183922 104802 183978
rect 104858 183922 104928 183978
rect 104608 183888 104928 183922
rect 135328 184350 135648 184384
rect 135328 184294 135398 184350
rect 135454 184294 135522 184350
rect 135578 184294 135648 184350
rect 135328 184226 135648 184294
rect 135328 184170 135398 184226
rect 135454 184170 135522 184226
rect 135578 184170 135648 184226
rect 135328 184102 135648 184170
rect 135328 184046 135398 184102
rect 135454 184046 135522 184102
rect 135578 184046 135648 184102
rect 135328 183978 135648 184046
rect 135328 183922 135398 183978
rect 135454 183922 135522 183978
rect 135578 183922 135648 183978
rect 135328 183888 135648 183922
rect 166048 184350 166368 184384
rect 166048 184294 166118 184350
rect 166174 184294 166242 184350
rect 166298 184294 166368 184350
rect 166048 184226 166368 184294
rect 166048 184170 166118 184226
rect 166174 184170 166242 184226
rect 166298 184170 166368 184226
rect 166048 184102 166368 184170
rect 166048 184046 166118 184102
rect 166174 184046 166242 184102
rect 166298 184046 166368 184102
rect 166048 183978 166368 184046
rect 166048 183922 166118 183978
rect 166174 183922 166242 183978
rect 166298 183922 166368 183978
rect 166048 183888 166368 183922
rect 196768 184350 197088 184384
rect 196768 184294 196838 184350
rect 196894 184294 196962 184350
rect 197018 184294 197088 184350
rect 196768 184226 197088 184294
rect 196768 184170 196838 184226
rect 196894 184170 196962 184226
rect 197018 184170 197088 184226
rect 196768 184102 197088 184170
rect 196768 184046 196838 184102
rect 196894 184046 196962 184102
rect 197018 184046 197088 184102
rect 196768 183978 197088 184046
rect 196768 183922 196838 183978
rect 196894 183922 196962 183978
rect 197018 183922 197088 183978
rect 196768 183888 197088 183922
rect 227488 184350 227808 184384
rect 227488 184294 227558 184350
rect 227614 184294 227682 184350
rect 227738 184294 227808 184350
rect 227488 184226 227808 184294
rect 227488 184170 227558 184226
rect 227614 184170 227682 184226
rect 227738 184170 227808 184226
rect 227488 184102 227808 184170
rect 227488 184046 227558 184102
rect 227614 184046 227682 184102
rect 227738 184046 227808 184102
rect 227488 183978 227808 184046
rect 227488 183922 227558 183978
rect 227614 183922 227682 183978
rect 227738 183922 227808 183978
rect 227488 183888 227808 183922
rect 258208 184350 258528 184384
rect 258208 184294 258278 184350
rect 258334 184294 258402 184350
rect 258458 184294 258528 184350
rect 258208 184226 258528 184294
rect 258208 184170 258278 184226
rect 258334 184170 258402 184226
rect 258458 184170 258528 184226
rect 258208 184102 258528 184170
rect 258208 184046 258278 184102
rect 258334 184046 258402 184102
rect 258458 184046 258528 184102
rect 258208 183978 258528 184046
rect 258208 183922 258278 183978
rect 258334 183922 258402 183978
rect 258458 183922 258528 183978
rect 258208 183888 258528 183922
rect 288928 184350 289248 184384
rect 288928 184294 288998 184350
rect 289054 184294 289122 184350
rect 289178 184294 289248 184350
rect 288928 184226 289248 184294
rect 288928 184170 288998 184226
rect 289054 184170 289122 184226
rect 289178 184170 289248 184226
rect 288928 184102 289248 184170
rect 288928 184046 288998 184102
rect 289054 184046 289122 184102
rect 289178 184046 289248 184102
rect 288928 183978 289248 184046
rect 288928 183922 288998 183978
rect 289054 183922 289122 183978
rect 289178 183922 289248 183978
rect 288928 183888 289248 183922
rect 319648 184350 319968 184384
rect 319648 184294 319718 184350
rect 319774 184294 319842 184350
rect 319898 184294 319968 184350
rect 319648 184226 319968 184294
rect 319648 184170 319718 184226
rect 319774 184170 319842 184226
rect 319898 184170 319968 184226
rect 319648 184102 319968 184170
rect 319648 184046 319718 184102
rect 319774 184046 319842 184102
rect 319898 184046 319968 184102
rect 319648 183978 319968 184046
rect 319648 183922 319718 183978
rect 319774 183922 319842 183978
rect 319898 183922 319968 183978
rect 319648 183888 319968 183922
rect 350368 184350 350688 184384
rect 350368 184294 350438 184350
rect 350494 184294 350562 184350
rect 350618 184294 350688 184350
rect 350368 184226 350688 184294
rect 350368 184170 350438 184226
rect 350494 184170 350562 184226
rect 350618 184170 350688 184226
rect 350368 184102 350688 184170
rect 350368 184046 350438 184102
rect 350494 184046 350562 184102
rect 350618 184046 350688 184102
rect 350368 183978 350688 184046
rect 350368 183922 350438 183978
rect 350494 183922 350562 183978
rect 350618 183922 350688 183978
rect 350368 183888 350688 183922
rect 381088 184350 381408 184384
rect 381088 184294 381158 184350
rect 381214 184294 381282 184350
rect 381338 184294 381408 184350
rect 381088 184226 381408 184294
rect 381088 184170 381158 184226
rect 381214 184170 381282 184226
rect 381338 184170 381408 184226
rect 381088 184102 381408 184170
rect 381088 184046 381158 184102
rect 381214 184046 381282 184102
rect 381338 184046 381408 184102
rect 381088 183978 381408 184046
rect 381088 183922 381158 183978
rect 381214 183922 381282 183978
rect 381338 183922 381408 183978
rect 381088 183888 381408 183922
rect 411808 184350 412128 184384
rect 411808 184294 411878 184350
rect 411934 184294 412002 184350
rect 412058 184294 412128 184350
rect 411808 184226 412128 184294
rect 411808 184170 411878 184226
rect 411934 184170 412002 184226
rect 412058 184170 412128 184226
rect 411808 184102 412128 184170
rect 411808 184046 411878 184102
rect 411934 184046 412002 184102
rect 412058 184046 412128 184102
rect 411808 183978 412128 184046
rect 411808 183922 411878 183978
rect 411934 183922 412002 183978
rect 412058 183922 412128 183978
rect 411808 183888 412128 183922
rect 442528 184350 442848 184384
rect 442528 184294 442598 184350
rect 442654 184294 442722 184350
rect 442778 184294 442848 184350
rect 442528 184226 442848 184294
rect 442528 184170 442598 184226
rect 442654 184170 442722 184226
rect 442778 184170 442848 184226
rect 442528 184102 442848 184170
rect 442528 184046 442598 184102
rect 442654 184046 442722 184102
rect 442778 184046 442848 184102
rect 442528 183978 442848 184046
rect 442528 183922 442598 183978
rect 442654 183922 442722 183978
rect 442778 183922 442848 183978
rect 442528 183888 442848 183922
rect 473248 184350 473568 184384
rect 473248 184294 473318 184350
rect 473374 184294 473442 184350
rect 473498 184294 473568 184350
rect 473248 184226 473568 184294
rect 473248 184170 473318 184226
rect 473374 184170 473442 184226
rect 473498 184170 473568 184226
rect 473248 184102 473568 184170
rect 473248 184046 473318 184102
rect 473374 184046 473442 184102
rect 473498 184046 473568 184102
rect 473248 183978 473568 184046
rect 473248 183922 473318 183978
rect 473374 183922 473442 183978
rect 473498 183922 473568 183978
rect 473248 183888 473568 183922
rect 503968 184350 504288 184384
rect 503968 184294 504038 184350
rect 504094 184294 504162 184350
rect 504218 184294 504288 184350
rect 503968 184226 504288 184294
rect 503968 184170 504038 184226
rect 504094 184170 504162 184226
rect 504218 184170 504288 184226
rect 503968 184102 504288 184170
rect 503968 184046 504038 184102
rect 504094 184046 504162 184102
rect 504218 184046 504288 184102
rect 503968 183978 504288 184046
rect 503968 183922 504038 183978
rect 504094 183922 504162 183978
rect 504218 183922 504288 183978
rect 503968 183888 504288 183922
rect 534688 184350 535008 184384
rect 534688 184294 534758 184350
rect 534814 184294 534882 184350
rect 534938 184294 535008 184350
rect 534688 184226 535008 184294
rect 534688 184170 534758 184226
rect 534814 184170 534882 184226
rect 534938 184170 535008 184226
rect 534688 184102 535008 184170
rect 534688 184046 534758 184102
rect 534814 184046 534882 184102
rect 534938 184046 535008 184102
rect 534688 183978 535008 184046
rect 534688 183922 534758 183978
rect 534814 183922 534882 183978
rect 534938 183922 535008 183978
rect 534688 183888 535008 183922
rect 565408 184350 565728 184384
rect 565408 184294 565478 184350
rect 565534 184294 565602 184350
rect 565658 184294 565728 184350
rect 565408 184226 565728 184294
rect 565408 184170 565478 184226
rect 565534 184170 565602 184226
rect 565658 184170 565728 184226
rect 565408 184102 565728 184170
rect 565408 184046 565478 184102
rect 565534 184046 565602 184102
rect 565658 184046 565728 184102
rect 565408 183978 565728 184046
rect 565408 183922 565478 183978
rect 565534 183922 565602 183978
rect 565658 183922 565728 183978
rect 565408 183888 565728 183922
rect 585564 178500 585620 205324
rect 585676 200004 585732 231868
rect 587132 221508 587188 258188
rect 587132 221442 587188 221452
rect 589098 256350 589718 273922
rect 590492 297892 590548 297902
rect 590492 264516 590548 297836
rect 590492 264450 590548 264460
rect 592818 280350 593438 297922
rect 592818 280294 592914 280350
rect 592970 280294 593038 280350
rect 593094 280294 593162 280350
rect 593218 280294 593286 280350
rect 593342 280294 593438 280350
rect 592818 280226 593438 280294
rect 592818 280170 592914 280226
rect 592970 280170 593038 280226
rect 593094 280170 593162 280226
rect 593218 280170 593286 280226
rect 593342 280170 593438 280226
rect 592818 280102 593438 280170
rect 592818 280046 592914 280102
rect 592970 280046 593038 280102
rect 593094 280046 593162 280102
rect 593218 280046 593286 280102
rect 593342 280046 593438 280102
rect 592818 279978 593438 280046
rect 592818 279922 592914 279978
rect 592970 279922 593038 279978
rect 593094 279922 593162 279978
rect 593218 279922 593286 279978
rect 593342 279922 593438 279978
rect 589098 256294 589194 256350
rect 589250 256294 589318 256350
rect 589374 256294 589442 256350
rect 589498 256294 589566 256350
rect 589622 256294 589718 256350
rect 589098 256226 589718 256294
rect 589098 256170 589194 256226
rect 589250 256170 589318 256226
rect 589374 256170 589442 256226
rect 589498 256170 589566 256226
rect 589622 256170 589718 256226
rect 589098 256102 589718 256170
rect 589098 256046 589194 256102
rect 589250 256046 589318 256102
rect 589374 256046 589442 256102
rect 589498 256046 589566 256102
rect 589622 256046 589718 256102
rect 589098 255978 589718 256046
rect 589098 255922 589194 255978
rect 589250 255922 589318 255978
rect 589374 255922 589442 255978
rect 589498 255922 589566 255978
rect 589622 255922 589718 255978
rect 589098 238350 589718 255922
rect 592818 262350 593438 279922
rect 592818 262294 592914 262350
rect 592970 262294 593038 262350
rect 593094 262294 593162 262350
rect 593218 262294 593286 262350
rect 593342 262294 593438 262350
rect 592818 262226 593438 262294
rect 592818 262170 592914 262226
rect 592970 262170 593038 262226
rect 593094 262170 593162 262226
rect 593218 262170 593286 262226
rect 593342 262170 593438 262226
rect 592818 262102 593438 262170
rect 592818 262046 592914 262102
rect 592970 262046 593038 262102
rect 593094 262046 593162 262102
rect 593218 262046 593286 262102
rect 593342 262046 593438 262102
rect 592818 261978 593438 262046
rect 592818 261922 592914 261978
rect 592970 261922 593038 261978
rect 593094 261922 593162 261978
rect 593218 261922 593286 261978
rect 593342 261922 593438 261978
rect 589098 238294 589194 238350
rect 589250 238294 589318 238350
rect 589374 238294 589442 238350
rect 589498 238294 589566 238350
rect 589622 238294 589718 238350
rect 589098 238226 589718 238294
rect 589098 238170 589194 238226
rect 589250 238170 589318 238226
rect 589374 238170 589442 238226
rect 589498 238170 589566 238226
rect 589622 238170 589718 238226
rect 589098 238102 589718 238170
rect 589098 238046 589194 238102
rect 589250 238046 589318 238102
rect 589374 238046 589442 238102
rect 589498 238046 589566 238102
rect 589622 238046 589718 238102
rect 589098 237978 589718 238046
rect 589098 237922 589194 237978
rect 589250 237922 589318 237978
rect 589374 237922 589442 237978
rect 589498 237922 589566 237978
rect 589622 237922 589718 237978
rect 585676 199938 585732 199948
rect 589098 220350 589718 237922
rect 589098 220294 589194 220350
rect 589250 220294 589318 220350
rect 589374 220294 589442 220350
rect 589498 220294 589566 220350
rect 589622 220294 589718 220350
rect 589098 220226 589718 220294
rect 589098 220170 589194 220226
rect 589250 220170 589318 220226
rect 589374 220170 589442 220226
rect 589498 220170 589566 220226
rect 589622 220170 589718 220226
rect 589098 220102 589718 220170
rect 589098 220046 589194 220102
rect 589250 220046 589318 220102
rect 589374 220046 589442 220102
rect 589498 220046 589566 220102
rect 589622 220046 589718 220102
rect 589098 219978 589718 220046
rect 589098 219922 589194 219978
rect 589250 219922 589318 219978
rect 589374 219922 589442 219978
rect 589498 219922 589566 219978
rect 589622 219922 589718 219978
rect 589098 202350 589718 219922
rect 590492 245028 590548 245038
rect 590492 210756 590548 244972
rect 590492 210690 590548 210700
rect 592818 244350 593438 261922
rect 592818 244294 592914 244350
rect 592970 244294 593038 244350
rect 593094 244294 593162 244350
rect 593218 244294 593286 244350
rect 593342 244294 593438 244350
rect 592818 244226 593438 244294
rect 592818 244170 592914 244226
rect 592970 244170 593038 244226
rect 593094 244170 593162 244226
rect 593218 244170 593286 244226
rect 593342 244170 593438 244226
rect 592818 244102 593438 244170
rect 592818 244046 592914 244102
rect 592970 244046 593038 244102
rect 593094 244046 593162 244102
rect 593218 244046 593286 244102
rect 593342 244046 593438 244102
rect 592818 243978 593438 244046
rect 592818 243922 592914 243978
rect 592970 243922 593038 243978
rect 593094 243922 593162 243978
rect 593218 243922 593286 243978
rect 593342 243922 593438 243978
rect 592818 226350 593438 243922
rect 592818 226294 592914 226350
rect 592970 226294 593038 226350
rect 593094 226294 593162 226350
rect 593218 226294 593286 226350
rect 593342 226294 593438 226350
rect 592818 226226 593438 226294
rect 592818 226170 592914 226226
rect 592970 226170 593038 226226
rect 593094 226170 593162 226226
rect 593218 226170 593286 226226
rect 593342 226170 593438 226226
rect 592818 226102 593438 226170
rect 592818 226046 592914 226102
rect 592970 226046 593038 226102
rect 593094 226046 593162 226102
rect 593218 226046 593286 226102
rect 593342 226046 593438 226102
rect 592818 225978 593438 226046
rect 592818 225922 592914 225978
rect 592970 225922 593038 225978
rect 593094 225922 593162 225978
rect 593218 225922 593286 225978
rect 593342 225922 593438 225978
rect 589098 202294 589194 202350
rect 589250 202294 589318 202350
rect 589374 202294 589442 202350
rect 589498 202294 589566 202350
rect 589622 202294 589718 202350
rect 589098 202226 589718 202294
rect 589098 202170 589194 202226
rect 589250 202170 589318 202226
rect 589374 202170 589442 202226
rect 589498 202170 589566 202226
rect 589622 202170 589718 202226
rect 589098 202102 589718 202170
rect 589098 202046 589194 202102
rect 589250 202046 589318 202102
rect 589374 202046 589442 202102
rect 589498 202046 589566 202102
rect 589622 202046 589718 202102
rect 589098 201978 589718 202046
rect 589098 201922 589194 201978
rect 589250 201922 589318 201978
rect 589374 201922 589442 201978
rect 589498 201922 589566 201978
rect 589622 201922 589718 201978
rect 585564 178434 585620 178444
rect 585676 192164 585732 192174
rect 27808 172350 28128 172384
rect 27808 172294 27878 172350
rect 27934 172294 28002 172350
rect 28058 172294 28128 172350
rect 27808 172226 28128 172294
rect 27808 172170 27878 172226
rect 27934 172170 28002 172226
rect 28058 172170 28128 172226
rect 27808 172102 28128 172170
rect 27808 172046 27878 172102
rect 27934 172046 28002 172102
rect 28058 172046 28128 172102
rect 27808 171978 28128 172046
rect 27808 171922 27878 171978
rect 27934 171922 28002 171978
rect 28058 171922 28128 171978
rect 27808 171888 28128 171922
rect 58528 172350 58848 172384
rect 58528 172294 58598 172350
rect 58654 172294 58722 172350
rect 58778 172294 58848 172350
rect 58528 172226 58848 172294
rect 58528 172170 58598 172226
rect 58654 172170 58722 172226
rect 58778 172170 58848 172226
rect 58528 172102 58848 172170
rect 58528 172046 58598 172102
rect 58654 172046 58722 172102
rect 58778 172046 58848 172102
rect 58528 171978 58848 172046
rect 58528 171922 58598 171978
rect 58654 171922 58722 171978
rect 58778 171922 58848 171978
rect 58528 171888 58848 171922
rect 89248 172350 89568 172384
rect 89248 172294 89318 172350
rect 89374 172294 89442 172350
rect 89498 172294 89568 172350
rect 89248 172226 89568 172294
rect 89248 172170 89318 172226
rect 89374 172170 89442 172226
rect 89498 172170 89568 172226
rect 89248 172102 89568 172170
rect 89248 172046 89318 172102
rect 89374 172046 89442 172102
rect 89498 172046 89568 172102
rect 89248 171978 89568 172046
rect 89248 171922 89318 171978
rect 89374 171922 89442 171978
rect 89498 171922 89568 171978
rect 89248 171888 89568 171922
rect 119968 172350 120288 172384
rect 119968 172294 120038 172350
rect 120094 172294 120162 172350
rect 120218 172294 120288 172350
rect 119968 172226 120288 172294
rect 119968 172170 120038 172226
rect 120094 172170 120162 172226
rect 120218 172170 120288 172226
rect 119968 172102 120288 172170
rect 119968 172046 120038 172102
rect 120094 172046 120162 172102
rect 120218 172046 120288 172102
rect 119968 171978 120288 172046
rect 119968 171922 120038 171978
rect 120094 171922 120162 171978
rect 120218 171922 120288 171978
rect 119968 171888 120288 171922
rect 150688 172350 151008 172384
rect 150688 172294 150758 172350
rect 150814 172294 150882 172350
rect 150938 172294 151008 172350
rect 150688 172226 151008 172294
rect 150688 172170 150758 172226
rect 150814 172170 150882 172226
rect 150938 172170 151008 172226
rect 150688 172102 151008 172170
rect 150688 172046 150758 172102
rect 150814 172046 150882 172102
rect 150938 172046 151008 172102
rect 150688 171978 151008 172046
rect 150688 171922 150758 171978
rect 150814 171922 150882 171978
rect 150938 171922 151008 171978
rect 150688 171888 151008 171922
rect 181408 172350 181728 172384
rect 181408 172294 181478 172350
rect 181534 172294 181602 172350
rect 181658 172294 181728 172350
rect 181408 172226 181728 172294
rect 181408 172170 181478 172226
rect 181534 172170 181602 172226
rect 181658 172170 181728 172226
rect 181408 172102 181728 172170
rect 181408 172046 181478 172102
rect 181534 172046 181602 172102
rect 181658 172046 181728 172102
rect 181408 171978 181728 172046
rect 181408 171922 181478 171978
rect 181534 171922 181602 171978
rect 181658 171922 181728 171978
rect 181408 171888 181728 171922
rect 212128 172350 212448 172384
rect 212128 172294 212198 172350
rect 212254 172294 212322 172350
rect 212378 172294 212448 172350
rect 212128 172226 212448 172294
rect 212128 172170 212198 172226
rect 212254 172170 212322 172226
rect 212378 172170 212448 172226
rect 212128 172102 212448 172170
rect 212128 172046 212198 172102
rect 212254 172046 212322 172102
rect 212378 172046 212448 172102
rect 212128 171978 212448 172046
rect 212128 171922 212198 171978
rect 212254 171922 212322 171978
rect 212378 171922 212448 171978
rect 212128 171888 212448 171922
rect 242848 172350 243168 172384
rect 242848 172294 242918 172350
rect 242974 172294 243042 172350
rect 243098 172294 243168 172350
rect 242848 172226 243168 172294
rect 242848 172170 242918 172226
rect 242974 172170 243042 172226
rect 243098 172170 243168 172226
rect 242848 172102 243168 172170
rect 242848 172046 242918 172102
rect 242974 172046 243042 172102
rect 243098 172046 243168 172102
rect 242848 171978 243168 172046
rect 242848 171922 242918 171978
rect 242974 171922 243042 171978
rect 243098 171922 243168 171978
rect 242848 171888 243168 171922
rect 273568 172350 273888 172384
rect 273568 172294 273638 172350
rect 273694 172294 273762 172350
rect 273818 172294 273888 172350
rect 273568 172226 273888 172294
rect 273568 172170 273638 172226
rect 273694 172170 273762 172226
rect 273818 172170 273888 172226
rect 273568 172102 273888 172170
rect 273568 172046 273638 172102
rect 273694 172046 273762 172102
rect 273818 172046 273888 172102
rect 273568 171978 273888 172046
rect 273568 171922 273638 171978
rect 273694 171922 273762 171978
rect 273818 171922 273888 171978
rect 273568 171888 273888 171922
rect 304288 172350 304608 172384
rect 304288 172294 304358 172350
rect 304414 172294 304482 172350
rect 304538 172294 304608 172350
rect 304288 172226 304608 172294
rect 304288 172170 304358 172226
rect 304414 172170 304482 172226
rect 304538 172170 304608 172226
rect 304288 172102 304608 172170
rect 304288 172046 304358 172102
rect 304414 172046 304482 172102
rect 304538 172046 304608 172102
rect 304288 171978 304608 172046
rect 304288 171922 304358 171978
rect 304414 171922 304482 171978
rect 304538 171922 304608 171978
rect 304288 171888 304608 171922
rect 335008 172350 335328 172384
rect 335008 172294 335078 172350
rect 335134 172294 335202 172350
rect 335258 172294 335328 172350
rect 335008 172226 335328 172294
rect 335008 172170 335078 172226
rect 335134 172170 335202 172226
rect 335258 172170 335328 172226
rect 335008 172102 335328 172170
rect 335008 172046 335078 172102
rect 335134 172046 335202 172102
rect 335258 172046 335328 172102
rect 335008 171978 335328 172046
rect 335008 171922 335078 171978
rect 335134 171922 335202 171978
rect 335258 171922 335328 171978
rect 335008 171888 335328 171922
rect 365728 172350 366048 172384
rect 365728 172294 365798 172350
rect 365854 172294 365922 172350
rect 365978 172294 366048 172350
rect 365728 172226 366048 172294
rect 365728 172170 365798 172226
rect 365854 172170 365922 172226
rect 365978 172170 366048 172226
rect 365728 172102 366048 172170
rect 365728 172046 365798 172102
rect 365854 172046 365922 172102
rect 365978 172046 366048 172102
rect 365728 171978 366048 172046
rect 365728 171922 365798 171978
rect 365854 171922 365922 171978
rect 365978 171922 366048 171978
rect 365728 171888 366048 171922
rect 396448 172350 396768 172384
rect 396448 172294 396518 172350
rect 396574 172294 396642 172350
rect 396698 172294 396768 172350
rect 396448 172226 396768 172294
rect 396448 172170 396518 172226
rect 396574 172170 396642 172226
rect 396698 172170 396768 172226
rect 396448 172102 396768 172170
rect 396448 172046 396518 172102
rect 396574 172046 396642 172102
rect 396698 172046 396768 172102
rect 396448 171978 396768 172046
rect 396448 171922 396518 171978
rect 396574 171922 396642 171978
rect 396698 171922 396768 171978
rect 396448 171888 396768 171922
rect 427168 172350 427488 172384
rect 427168 172294 427238 172350
rect 427294 172294 427362 172350
rect 427418 172294 427488 172350
rect 427168 172226 427488 172294
rect 427168 172170 427238 172226
rect 427294 172170 427362 172226
rect 427418 172170 427488 172226
rect 427168 172102 427488 172170
rect 427168 172046 427238 172102
rect 427294 172046 427362 172102
rect 427418 172046 427488 172102
rect 427168 171978 427488 172046
rect 427168 171922 427238 171978
rect 427294 171922 427362 171978
rect 427418 171922 427488 171978
rect 427168 171888 427488 171922
rect 457888 172350 458208 172384
rect 457888 172294 457958 172350
rect 458014 172294 458082 172350
rect 458138 172294 458208 172350
rect 457888 172226 458208 172294
rect 457888 172170 457958 172226
rect 458014 172170 458082 172226
rect 458138 172170 458208 172226
rect 457888 172102 458208 172170
rect 457888 172046 457958 172102
rect 458014 172046 458082 172102
rect 458138 172046 458208 172102
rect 457888 171978 458208 172046
rect 457888 171922 457958 171978
rect 458014 171922 458082 171978
rect 458138 171922 458208 171978
rect 457888 171888 458208 171922
rect 488608 172350 488928 172384
rect 488608 172294 488678 172350
rect 488734 172294 488802 172350
rect 488858 172294 488928 172350
rect 488608 172226 488928 172294
rect 488608 172170 488678 172226
rect 488734 172170 488802 172226
rect 488858 172170 488928 172226
rect 488608 172102 488928 172170
rect 488608 172046 488678 172102
rect 488734 172046 488802 172102
rect 488858 172046 488928 172102
rect 488608 171978 488928 172046
rect 488608 171922 488678 171978
rect 488734 171922 488802 171978
rect 488858 171922 488928 171978
rect 488608 171888 488928 171922
rect 519328 172350 519648 172384
rect 519328 172294 519398 172350
rect 519454 172294 519522 172350
rect 519578 172294 519648 172350
rect 519328 172226 519648 172294
rect 519328 172170 519398 172226
rect 519454 172170 519522 172226
rect 519578 172170 519648 172226
rect 519328 172102 519648 172170
rect 519328 172046 519398 172102
rect 519454 172046 519522 172102
rect 519578 172046 519648 172102
rect 519328 171978 519648 172046
rect 519328 171922 519398 171978
rect 519454 171922 519522 171978
rect 519578 171922 519648 171978
rect 519328 171888 519648 171922
rect 550048 172350 550368 172384
rect 550048 172294 550118 172350
rect 550174 172294 550242 172350
rect 550298 172294 550368 172350
rect 550048 172226 550368 172294
rect 550048 172170 550118 172226
rect 550174 172170 550242 172226
rect 550298 172170 550368 172226
rect 550048 172102 550368 172170
rect 550048 172046 550118 172102
rect 550174 172046 550242 172102
rect 550298 172046 550368 172102
rect 550048 171978 550368 172046
rect 550048 171922 550118 171978
rect 550174 171922 550242 171978
rect 550298 171922 550368 171978
rect 550048 171888 550368 171922
rect 585676 167748 585732 192108
rect 589098 184350 589718 201922
rect 589098 184294 589194 184350
rect 589250 184294 589318 184350
rect 589374 184294 589442 184350
rect 589498 184294 589566 184350
rect 589622 184294 589718 184350
rect 589098 184226 589718 184294
rect 589098 184170 589194 184226
rect 589250 184170 589318 184226
rect 589374 184170 589442 184226
rect 589498 184170 589566 184226
rect 589622 184170 589718 184226
rect 589098 184102 589718 184170
rect 589098 184046 589194 184102
rect 589250 184046 589318 184102
rect 589374 184046 589442 184102
rect 589498 184046 589566 184102
rect 589622 184046 589718 184102
rect 589098 183978 589718 184046
rect 589098 183922 589194 183978
rect 589250 183922 589318 183978
rect 589374 183922 589442 183978
rect 589498 183922 589566 183978
rect 589622 183922 589718 183978
rect 585676 167682 585732 167692
rect 585788 178948 585844 178958
rect 5418 166294 5514 166350
rect 5570 166294 5638 166350
rect 5694 166294 5762 166350
rect 5818 166294 5886 166350
rect 5942 166294 6038 166350
rect 5418 166226 6038 166294
rect 5418 166170 5514 166226
rect 5570 166170 5638 166226
rect 5694 166170 5762 166226
rect 5818 166170 5886 166226
rect 5942 166170 6038 166226
rect 5418 166102 6038 166170
rect 5418 166046 5514 166102
rect 5570 166046 5638 166102
rect 5694 166046 5762 166102
rect 5818 166046 5886 166102
rect 5942 166046 6038 166102
rect 5418 165978 6038 166046
rect 5418 165922 5514 165978
rect 5570 165922 5638 165978
rect 5694 165922 5762 165978
rect 5818 165922 5886 165978
rect 5942 165922 6038 165978
rect -956 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 -336 148350
rect -956 148226 -336 148294
rect -956 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 -336 148226
rect -956 148102 -336 148170
rect -956 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 -336 148102
rect -956 147978 -336 148046
rect -956 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 -336 147978
rect -956 130350 -336 147922
rect 4172 149716 4228 149726
rect 4172 133476 4228 149660
rect 5418 148350 6038 165922
rect 12448 166350 12768 166384
rect 12448 166294 12518 166350
rect 12574 166294 12642 166350
rect 12698 166294 12768 166350
rect 12448 166226 12768 166294
rect 12448 166170 12518 166226
rect 12574 166170 12642 166226
rect 12698 166170 12768 166226
rect 12448 166102 12768 166170
rect 12448 166046 12518 166102
rect 12574 166046 12642 166102
rect 12698 166046 12768 166102
rect 12448 165978 12768 166046
rect 12448 165922 12518 165978
rect 12574 165922 12642 165978
rect 12698 165922 12768 165978
rect 12448 165888 12768 165922
rect 43168 166350 43488 166384
rect 43168 166294 43238 166350
rect 43294 166294 43362 166350
rect 43418 166294 43488 166350
rect 43168 166226 43488 166294
rect 43168 166170 43238 166226
rect 43294 166170 43362 166226
rect 43418 166170 43488 166226
rect 43168 166102 43488 166170
rect 43168 166046 43238 166102
rect 43294 166046 43362 166102
rect 43418 166046 43488 166102
rect 43168 165978 43488 166046
rect 43168 165922 43238 165978
rect 43294 165922 43362 165978
rect 43418 165922 43488 165978
rect 43168 165888 43488 165922
rect 73888 166350 74208 166384
rect 73888 166294 73958 166350
rect 74014 166294 74082 166350
rect 74138 166294 74208 166350
rect 73888 166226 74208 166294
rect 73888 166170 73958 166226
rect 74014 166170 74082 166226
rect 74138 166170 74208 166226
rect 73888 166102 74208 166170
rect 73888 166046 73958 166102
rect 74014 166046 74082 166102
rect 74138 166046 74208 166102
rect 73888 165978 74208 166046
rect 73888 165922 73958 165978
rect 74014 165922 74082 165978
rect 74138 165922 74208 165978
rect 73888 165888 74208 165922
rect 104608 166350 104928 166384
rect 104608 166294 104678 166350
rect 104734 166294 104802 166350
rect 104858 166294 104928 166350
rect 104608 166226 104928 166294
rect 104608 166170 104678 166226
rect 104734 166170 104802 166226
rect 104858 166170 104928 166226
rect 104608 166102 104928 166170
rect 104608 166046 104678 166102
rect 104734 166046 104802 166102
rect 104858 166046 104928 166102
rect 104608 165978 104928 166046
rect 104608 165922 104678 165978
rect 104734 165922 104802 165978
rect 104858 165922 104928 165978
rect 104608 165888 104928 165922
rect 135328 166350 135648 166384
rect 135328 166294 135398 166350
rect 135454 166294 135522 166350
rect 135578 166294 135648 166350
rect 135328 166226 135648 166294
rect 135328 166170 135398 166226
rect 135454 166170 135522 166226
rect 135578 166170 135648 166226
rect 135328 166102 135648 166170
rect 135328 166046 135398 166102
rect 135454 166046 135522 166102
rect 135578 166046 135648 166102
rect 135328 165978 135648 166046
rect 135328 165922 135398 165978
rect 135454 165922 135522 165978
rect 135578 165922 135648 165978
rect 135328 165888 135648 165922
rect 166048 166350 166368 166384
rect 166048 166294 166118 166350
rect 166174 166294 166242 166350
rect 166298 166294 166368 166350
rect 166048 166226 166368 166294
rect 166048 166170 166118 166226
rect 166174 166170 166242 166226
rect 166298 166170 166368 166226
rect 166048 166102 166368 166170
rect 166048 166046 166118 166102
rect 166174 166046 166242 166102
rect 166298 166046 166368 166102
rect 166048 165978 166368 166046
rect 166048 165922 166118 165978
rect 166174 165922 166242 165978
rect 166298 165922 166368 165978
rect 166048 165888 166368 165922
rect 196768 166350 197088 166384
rect 196768 166294 196838 166350
rect 196894 166294 196962 166350
rect 197018 166294 197088 166350
rect 196768 166226 197088 166294
rect 196768 166170 196838 166226
rect 196894 166170 196962 166226
rect 197018 166170 197088 166226
rect 196768 166102 197088 166170
rect 196768 166046 196838 166102
rect 196894 166046 196962 166102
rect 197018 166046 197088 166102
rect 196768 165978 197088 166046
rect 196768 165922 196838 165978
rect 196894 165922 196962 165978
rect 197018 165922 197088 165978
rect 196768 165888 197088 165922
rect 227488 166350 227808 166384
rect 227488 166294 227558 166350
rect 227614 166294 227682 166350
rect 227738 166294 227808 166350
rect 227488 166226 227808 166294
rect 227488 166170 227558 166226
rect 227614 166170 227682 166226
rect 227738 166170 227808 166226
rect 227488 166102 227808 166170
rect 227488 166046 227558 166102
rect 227614 166046 227682 166102
rect 227738 166046 227808 166102
rect 227488 165978 227808 166046
rect 227488 165922 227558 165978
rect 227614 165922 227682 165978
rect 227738 165922 227808 165978
rect 227488 165888 227808 165922
rect 258208 166350 258528 166384
rect 258208 166294 258278 166350
rect 258334 166294 258402 166350
rect 258458 166294 258528 166350
rect 258208 166226 258528 166294
rect 258208 166170 258278 166226
rect 258334 166170 258402 166226
rect 258458 166170 258528 166226
rect 258208 166102 258528 166170
rect 258208 166046 258278 166102
rect 258334 166046 258402 166102
rect 258458 166046 258528 166102
rect 258208 165978 258528 166046
rect 258208 165922 258278 165978
rect 258334 165922 258402 165978
rect 258458 165922 258528 165978
rect 258208 165888 258528 165922
rect 288928 166350 289248 166384
rect 288928 166294 288998 166350
rect 289054 166294 289122 166350
rect 289178 166294 289248 166350
rect 288928 166226 289248 166294
rect 288928 166170 288998 166226
rect 289054 166170 289122 166226
rect 289178 166170 289248 166226
rect 288928 166102 289248 166170
rect 288928 166046 288998 166102
rect 289054 166046 289122 166102
rect 289178 166046 289248 166102
rect 288928 165978 289248 166046
rect 288928 165922 288998 165978
rect 289054 165922 289122 165978
rect 289178 165922 289248 165978
rect 288928 165888 289248 165922
rect 319648 166350 319968 166384
rect 319648 166294 319718 166350
rect 319774 166294 319842 166350
rect 319898 166294 319968 166350
rect 319648 166226 319968 166294
rect 319648 166170 319718 166226
rect 319774 166170 319842 166226
rect 319898 166170 319968 166226
rect 319648 166102 319968 166170
rect 319648 166046 319718 166102
rect 319774 166046 319842 166102
rect 319898 166046 319968 166102
rect 319648 165978 319968 166046
rect 319648 165922 319718 165978
rect 319774 165922 319842 165978
rect 319898 165922 319968 165978
rect 319648 165888 319968 165922
rect 350368 166350 350688 166384
rect 350368 166294 350438 166350
rect 350494 166294 350562 166350
rect 350618 166294 350688 166350
rect 350368 166226 350688 166294
rect 350368 166170 350438 166226
rect 350494 166170 350562 166226
rect 350618 166170 350688 166226
rect 350368 166102 350688 166170
rect 350368 166046 350438 166102
rect 350494 166046 350562 166102
rect 350618 166046 350688 166102
rect 350368 165978 350688 166046
rect 350368 165922 350438 165978
rect 350494 165922 350562 165978
rect 350618 165922 350688 165978
rect 350368 165888 350688 165922
rect 381088 166350 381408 166384
rect 381088 166294 381158 166350
rect 381214 166294 381282 166350
rect 381338 166294 381408 166350
rect 381088 166226 381408 166294
rect 381088 166170 381158 166226
rect 381214 166170 381282 166226
rect 381338 166170 381408 166226
rect 381088 166102 381408 166170
rect 381088 166046 381158 166102
rect 381214 166046 381282 166102
rect 381338 166046 381408 166102
rect 381088 165978 381408 166046
rect 381088 165922 381158 165978
rect 381214 165922 381282 165978
rect 381338 165922 381408 165978
rect 381088 165888 381408 165922
rect 411808 166350 412128 166384
rect 411808 166294 411878 166350
rect 411934 166294 412002 166350
rect 412058 166294 412128 166350
rect 411808 166226 412128 166294
rect 411808 166170 411878 166226
rect 411934 166170 412002 166226
rect 412058 166170 412128 166226
rect 411808 166102 412128 166170
rect 411808 166046 411878 166102
rect 411934 166046 412002 166102
rect 412058 166046 412128 166102
rect 411808 165978 412128 166046
rect 411808 165922 411878 165978
rect 411934 165922 412002 165978
rect 412058 165922 412128 165978
rect 411808 165888 412128 165922
rect 442528 166350 442848 166384
rect 442528 166294 442598 166350
rect 442654 166294 442722 166350
rect 442778 166294 442848 166350
rect 442528 166226 442848 166294
rect 442528 166170 442598 166226
rect 442654 166170 442722 166226
rect 442778 166170 442848 166226
rect 442528 166102 442848 166170
rect 442528 166046 442598 166102
rect 442654 166046 442722 166102
rect 442778 166046 442848 166102
rect 442528 165978 442848 166046
rect 442528 165922 442598 165978
rect 442654 165922 442722 165978
rect 442778 165922 442848 165978
rect 442528 165888 442848 165922
rect 473248 166350 473568 166384
rect 473248 166294 473318 166350
rect 473374 166294 473442 166350
rect 473498 166294 473568 166350
rect 473248 166226 473568 166294
rect 473248 166170 473318 166226
rect 473374 166170 473442 166226
rect 473498 166170 473568 166226
rect 473248 166102 473568 166170
rect 473248 166046 473318 166102
rect 473374 166046 473442 166102
rect 473498 166046 473568 166102
rect 473248 165978 473568 166046
rect 473248 165922 473318 165978
rect 473374 165922 473442 165978
rect 473498 165922 473568 165978
rect 473248 165888 473568 165922
rect 503968 166350 504288 166384
rect 503968 166294 504038 166350
rect 504094 166294 504162 166350
rect 504218 166294 504288 166350
rect 503968 166226 504288 166294
rect 503968 166170 504038 166226
rect 504094 166170 504162 166226
rect 504218 166170 504288 166226
rect 503968 166102 504288 166170
rect 503968 166046 504038 166102
rect 504094 166046 504162 166102
rect 504218 166046 504288 166102
rect 503968 165978 504288 166046
rect 503968 165922 504038 165978
rect 504094 165922 504162 165978
rect 504218 165922 504288 165978
rect 503968 165888 504288 165922
rect 534688 166350 535008 166384
rect 534688 166294 534758 166350
rect 534814 166294 534882 166350
rect 534938 166294 535008 166350
rect 534688 166226 535008 166294
rect 534688 166170 534758 166226
rect 534814 166170 534882 166226
rect 534938 166170 535008 166226
rect 534688 166102 535008 166170
rect 534688 166046 534758 166102
rect 534814 166046 534882 166102
rect 534938 166046 535008 166102
rect 534688 165978 535008 166046
rect 534688 165922 534758 165978
rect 534814 165922 534882 165978
rect 534938 165922 535008 165978
rect 534688 165888 535008 165922
rect 565408 166350 565728 166384
rect 565408 166294 565478 166350
rect 565534 166294 565602 166350
rect 565658 166294 565728 166350
rect 565408 166226 565728 166294
rect 565408 166170 565478 166226
rect 565534 166170 565602 166226
rect 565658 166170 565728 166226
rect 565408 166102 565728 166170
rect 565408 166046 565478 166102
rect 565534 166046 565602 166102
rect 565658 166046 565728 166102
rect 565408 165978 565728 166046
rect 565408 165922 565478 165978
rect 565534 165922 565602 165978
rect 565658 165922 565728 165978
rect 565408 165888 565728 165922
rect 585452 165732 585508 165742
rect 5418 148294 5514 148350
rect 5570 148294 5638 148350
rect 5694 148294 5762 148350
rect 5818 148294 5886 148350
rect 5942 148294 6038 148350
rect 5418 148226 6038 148294
rect 5418 148170 5514 148226
rect 5570 148170 5638 148226
rect 5694 148170 5762 148226
rect 5818 148170 5886 148226
rect 5942 148170 6038 148226
rect 5418 148102 6038 148170
rect 5418 148046 5514 148102
rect 5570 148046 5638 148102
rect 5694 148046 5762 148102
rect 5818 148046 5886 148102
rect 5942 148046 6038 148102
rect 5418 147978 6038 148046
rect 5418 147922 5514 147978
rect 5570 147922 5638 147978
rect 5694 147922 5762 147978
rect 5818 147922 5886 147978
rect 5942 147922 6038 147978
rect 4172 133410 4228 133420
rect 4284 135604 4340 135614
rect -956 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 -336 130350
rect -956 130226 -336 130294
rect -956 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 -336 130226
rect -956 130102 -336 130170
rect -956 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 -336 130102
rect -956 129978 -336 130046
rect -956 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 -336 129978
rect -956 112350 -336 129922
rect 4284 122948 4340 135548
rect 4284 122882 4340 122892
rect 5418 130350 6038 147922
rect 6188 163828 6244 163838
rect 6188 144004 6244 163772
rect 27808 154350 28128 154384
rect 27808 154294 27878 154350
rect 27934 154294 28002 154350
rect 28058 154294 28128 154350
rect 27808 154226 28128 154294
rect 27808 154170 27878 154226
rect 27934 154170 28002 154226
rect 28058 154170 28128 154226
rect 27808 154102 28128 154170
rect 27808 154046 27878 154102
rect 27934 154046 28002 154102
rect 28058 154046 28128 154102
rect 27808 153978 28128 154046
rect 27808 153922 27878 153978
rect 27934 153922 28002 153978
rect 28058 153922 28128 153978
rect 27808 153888 28128 153922
rect 58528 154350 58848 154384
rect 58528 154294 58598 154350
rect 58654 154294 58722 154350
rect 58778 154294 58848 154350
rect 58528 154226 58848 154294
rect 58528 154170 58598 154226
rect 58654 154170 58722 154226
rect 58778 154170 58848 154226
rect 58528 154102 58848 154170
rect 58528 154046 58598 154102
rect 58654 154046 58722 154102
rect 58778 154046 58848 154102
rect 58528 153978 58848 154046
rect 58528 153922 58598 153978
rect 58654 153922 58722 153978
rect 58778 153922 58848 153978
rect 58528 153888 58848 153922
rect 89248 154350 89568 154384
rect 89248 154294 89318 154350
rect 89374 154294 89442 154350
rect 89498 154294 89568 154350
rect 89248 154226 89568 154294
rect 89248 154170 89318 154226
rect 89374 154170 89442 154226
rect 89498 154170 89568 154226
rect 89248 154102 89568 154170
rect 89248 154046 89318 154102
rect 89374 154046 89442 154102
rect 89498 154046 89568 154102
rect 89248 153978 89568 154046
rect 89248 153922 89318 153978
rect 89374 153922 89442 153978
rect 89498 153922 89568 153978
rect 89248 153888 89568 153922
rect 119968 154350 120288 154384
rect 119968 154294 120038 154350
rect 120094 154294 120162 154350
rect 120218 154294 120288 154350
rect 119968 154226 120288 154294
rect 119968 154170 120038 154226
rect 120094 154170 120162 154226
rect 120218 154170 120288 154226
rect 119968 154102 120288 154170
rect 119968 154046 120038 154102
rect 120094 154046 120162 154102
rect 120218 154046 120288 154102
rect 119968 153978 120288 154046
rect 119968 153922 120038 153978
rect 120094 153922 120162 153978
rect 120218 153922 120288 153978
rect 119968 153888 120288 153922
rect 150688 154350 151008 154384
rect 150688 154294 150758 154350
rect 150814 154294 150882 154350
rect 150938 154294 151008 154350
rect 150688 154226 151008 154294
rect 150688 154170 150758 154226
rect 150814 154170 150882 154226
rect 150938 154170 151008 154226
rect 150688 154102 151008 154170
rect 150688 154046 150758 154102
rect 150814 154046 150882 154102
rect 150938 154046 151008 154102
rect 150688 153978 151008 154046
rect 150688 153922 150758 153978
rect 150814 153922 150882 153978
rect 150938 153922 151008 153978
rect 150688 153888 151008 153922
rect 181408 154350 181728 154384
rect 181408 154294 181478 154350
rect 181534 154294 181602 154350
rect 181658 154294 181728 154350
rect 181408 154226 181728 154294
rect 181408 154170 181478 154226
rect 181534 154170 181602 154226
rect 181658 154170 181728 154226
rect 181408 154102 181728 154170
rect 181408 154046 181478 154102
rect 181534 154046 181602 154102
rect 181658 154046 181728 154102
rect 181408 153978 181728 154046
rect 181408 153922 181478 153978
rect 181534 153922 181602 153978
rect 181658 153922 181728 153978
rect 181408 153888 181728 153922
rect 212128 154350 212448 154384
rect 212128 154294 212198 154350
rect 212254 154294 212322 154350
rect 212378 154294 212448 154350
rect 212128 154226 212448 154294
rect 212128 154170 212198 154226
rect 212254 154170 212322 154226
rect 212378 154170 212448 154226
rect 212128 154102 212448 154170
rect 212128 154046 212198 154102
rect 212254 154046 212322 154102
rect 212378 154046 212448 154102
rect 212128 153978 212448 154046
rect 212128 153922 212198 153978
rect 212254 153922 212322 153978
rect 212378 153922 212448 153978
rect 212128 153888 212448 153922
rect 242848 154350 243168 154384
rect 242848 154294 242918 154350
rect 242974 154294 243042 154350
rect 243098 154294 243168 154350
rect 242848 154226 243168 154294
rect 242848 154170 242918 154226
rect 242974 154170 243042 154226
rect 243098 154170 243168 154226
rect 242848 154102 243168 154170
rect 242848 154046 242918 154102
rect 242974 154046 243042 154102
rect 243098 154046 243168 154102
rect 242848 153978 243168 154046
rect 242848 153922 242918 153978
rect 242974 153922 243042 153978
rect 243098 153922 243168 153978
rect 242848 153888 243168 153922
rect 273568 154350 273888 154384
rect 273568 154294 273638 154350
rect 273694 154294 273762 154350
rect 273818 154294 273888 154350
rect 273568 154226 273888 154294
rect 273568 154170 273638 154226
rect 273694 154170 273762 154226
rect 273818 154170 273888 154226
rect 273568 154102 273888 154170
rect 273568 154046 273638 154102
rect 273694 154046 273762 154102
rect 273818 154046 273888 154102
rect 273568 153978 273888 154046
rect 273568 153922 273638 153978
rect 273694 153922 273762 153978
rect 273818 153922 273888 153978
rect 273568 153888 273888 153922
rect 304288 154350 304608 154384
rect 304288 154294 304358 154350
rect 304414 154294 304482 154350
rect 304538 154294 304608 154350
rect 304288 154226 304608 154294
rect 304288 154170 304358 154226
rect 304414 154170 304482 154226
rect 304538 154170 304608 154226
rect 304288 154102 304608 154170
rect 304288 154046 304358 154102
rect 304414 154046 304482 154102
rect 304538 154046 304608 154102
rect 304288 153978 304608 154046
rect 304288 153922 304358 153978
rect 304414 153922 304482 153978
rect 304538 153922 304608 153978
rect 304288 153888 304608 153922
rect 335008 154350 335328 154384
rect 335008 154294 335078 154350
rect 335134 154294 335202 154350
rect 335258 154294 335328 154350
rect 335008 154226 335328 154294
rect 335008 154170 335078 154226
rect 335134 154170 335202 154226
rect 335258 154170 335328 154226
rect 335008 154102 335328 154170
rect 335008 154046 335078 154102
rect 335134 154046 335202 154102
rect 335258 154046 335328 154102
rect 335008 153978 335328 154046
rect 335008 153922 335078 153978
rect 335134 153922 335202 153978
rect 335258 153922 335328 153978
rect 335008 153888 335328 153922
rect 365728 154350 366048 154384
rect 365728 154294 365798 154350
rect 365854 154294 365922 154350
rect 365978 154294 366048 154350
rect 365728 154226 366048 154294
rect 365728 154170 365798 154226
rect 365854 154170 365922 154226
rect 365978 154170 366048 154226
rect 365728 154102 366048 154170
rect 365728 154046 365798 154102
rect 365854 154046 365922 154102
rect 365978 154046 366048 154102
rect 365728 153978 366048 154046
rect 365728 153922 365798 153978
rect 365854 153922 365922 153978
rect 365978 153922 366048 153978
rect 365728 153888 366048 153922
rect 396448 154350 396768 154384
rect 396448 154294 396518 154350
rect 396574 154294 396642 154350
rect 396698 154294 396768 154350
rect 396448 154226 396768 154294
rect 396448 154170 396518 154226
rect 396574 154170 396642 154226
rect 396698 154170 396768 154226
rect 396448 154102 396768 154170
rect 396448 154046 396518 154102
rect 396574 154046 396642 154102
rect 396698 154046 396768 154102
rect 396448 153978 396768 154046
rect 396448 153922 396518 153978
rect 396574 153922 396642 153978
rect 396698 153922 396768 153978
rect 396448 153888 396768 153922
rect 427168 154350 427488 154384
rect 427168 154294 427238 154350
rect 427294 154294 427362 154350
rect 427418 154294 427488 154350
rect 427168 154226 427488 154294
rect 427168 154170 427238 154226
rect 427294 154170 427362 154226
rect 427418 154170 427488 154226
rect 427168 154102 427488 154170
rect 427168 154046 427238 154102
rect 427294 154046 427362 154102
rect 427418 154046 427488 154102
rect 427168 153978 427488 154046
rect 427168 153922 427238 153978
rect 427294 153922 427362 153978
rect 427418 153922 427488 153978
rect 427168 153888 427488 153922
rect 457888 154350 458208 154384
rect 457888 154294 457958 154350
rect 458014 154294 458082 154350
rect 458138 154294 458208 154350
rect 457888 154226 458208 154294
rect 457888 154170 457958 154226
rect 458014 154170 458082 154226
rect 458138 154170 458208 154226
rect 457888 154102 458208 154170
rect 457888 154046 457958 154102
rect 458014 154046 458082 154102
rect 458138 154046 458208 154102
rect 457888 153978 458208 154046
rect 457888 153922 457958 153978
rect 458014 153922 458082 153978
rect 458138 153922 458208 153978
rect 457888 153888 458208 153922
rect 488608 154350 488928 154384
rect 488608 154294 488678 154350
rect 488734 154294 488802 154350
rect 488858 154294 488928 154350
rect 488608 154226 488928 154294
rect 488608 154170 488678 154226
rect 488734 154170 488802 154226
rect 488858 154170 488928 154226
rect 488608 154102 488928 154170
rect 488608 154046 488678 154102
rect 488734 154046 488802 154102
rect 488858 154046 488928 154102
rect 488608 153978 488928 154046
rect 488608 153922 488678 153978
rect 488734 153922 488802 153978
rect 488858 153922 488928 153978
rect 488608 153888 488928 153922
rect 519328 154350 519648 154384
rect 519328 154294 519398 154350
rect 519454 154294 519522 154350
rect 519578 154294 519648 154350
rect 519328 154226 519648 154294
rect 519328 154170 519398 154226
rect 519454 154170 519522 154226
rect 519578 154170 519648 154226
rect 519328 154102 519648 154170
rect 519328 154046 519398 154102
rect 519454 154046 519522 154102
rect 519578 154046 519648 154102
rect 519328 153978 519648 154046
rect 519328 153922 519398 153978
rect 519454 153922 519522 153978
rect 519578 153922 519648 153978
rect 519328 153888 519648 153922
rect 550048 154350 550368 154384
rect 550048 154294 550118 154350
rect 550174 154294 550242 154350
rect 550298 154294 550368 154350
rect 550048 154226 550368 154294
rect 550048 154170 550118 154226
rect 550174 154170 550242 154226
rect 550298 154170 550368 154226
rect 550048 154102 550368 154170
rect 550048 154046 550118 154102
rect 550174 154046 550242 154102
rect 550298 154046 550368 154102
rect 550048 153978 550368 154046
rect 550048 153922 550118 153978
rect 550174 153922 550242 153978
rect 550298 153922 550368 153978
rect 550048 153888 550368 153922
rect 12448 148350 12768 148384
rect 12448 148294 12518 148350
rect 12574 148294 12642 148350
rect 12698 148294 12768 148350
rect 12448 148226 12768 148294
rect 12448 148170 12518 148226
rect 12574 148170 12642 148226
rect 12698 148170 12768 148226
rect 12448 148102 12768 148170
rect 12448 148046 12518 148102
rect 12574 148046 12642 148102
rect 12698 148046 12768 148102
rect 12448 147978 12768 148046
rect 12448 147922 12518 147978
rect 12574 147922 12642 147978
rect 12698 147922 12768 147978
rect 12448 147888 12768 147922
rect 43168 148350 43488 148384
rect 43168 148294 43238 148350
rect 43294 148294 43362 148350
rect 43418 148294 43488 148350
rect 43168 148226 43488 148294
rect 43168 148170 43238 148226
rect 43294 148170 43362 148226
rect 43418 148170 43488 148226
rect 43168 148102 43488 148170
rect 43168 148046 43238 148102
rect 43294 148046 43362 148102
rect 43418 148046 43488 148102
rect 43168 147978 43488 148046
rect 43168 147922 43238 147978
rect 43294 147922 43362 147978
rect 43418 147922 43488 147978
rect 43168 147888 43488 147922
rect 73888 148350 74208 148384
rect 73888 148294 73958 148350
rect 74014 148294 74082 148350
rect 74138 148294 74208 148350
rect 73888 148226 74208 148294
rect 73888 148170 73958 148226
rect 74014 148170 74082 148226
rect 74138 148170 74208 148226
rect 73888 148102 74208 148170
rect 73888 148046 73958 148102
rect 74014 148046 74082 148102
rect 74138 148046 74208 148102
rect 73888 147978 74208 148046
rect 73888 147922 73958 147978
rect 74014 147922 74082 147978
rect 74138 147922 74208 147978
rect 73888 147888 74208 147922
rect 104608 148350 104928 148384
rect 104608 148294 104678 148350
rect 104734 148294 104802 148350
rect 104858 148294 104928 148350
rect 104608 148226 104928 148294
rect 104608 148170 104678 148226
rect 104734 148170 104802 148226
rect 104858 148170 104928 148226
rect 104608 148102 104928 148170
rect 104608 148046 104678 148102
rect 104734 148046 104802 148102
rect 104858 148046 104928 148102
rect 104608 147978 104928 148046
rect 104608 147922 104678 147978
rect 104734 147922 104802 147978
rect 104858 147922 104928 147978
rect 104608 147888 104928 147922
rect 135328 148350 135648 148384
rect 135328 148294 135398 148350
rect 135454 148294 135522 148350
rect 135578 148294 135648 148350
rect 135328 148226 135648 148294
rect 135328 148170 135398 148226
rect 135454 148170 135522 148226
rect 135578 148170 135648 148226
rect 135328 148102 135648 148170
rect 135328 148046 135398 148102
rect 135454 148046 135522 148102
rect 135578 148046 135648 148102
rect 135328 147978 135648 148046
rect 135328 147922 135398 147978
rect 135454 147922 135522 147978
rect 135578 147922 135648 147978
rect 135328 147888 135648 147922
rect 166048 148350 166368 148384
rect 166048 148294 166118 148350
rect 166174 148294 166242 148350
rect 166298 148294 166368 148350
rect 166048 148226 166368 148294
rect 166048 148170 166118 148226
rect 166174 148170 166242 148226
rect 166298 148170 166368 148226
rect 166048 148102 166368 148170
rect 166048 148046 166118 148102
rect 166174 148046 166242 148102
rect 166298 148046 166368 148102
rect 166048 147978 166368 148046
rect 166048 147922 166118 147978
rect 166174 147922 166242 147978
rect 166298 147922 166368 147978
rect 166048 147888 166368 147922
rect 196768 148350 197088 148384
rect 196768 148294 196838 148350
rect 196894 148294 196962 148350
rect 197018 148294 197088 148350
rect 196768 148226 197088 148294
rect 196768 148170 196838 148226
rect 196894 148170 196962 148226
rect 197018 148170 197088 148226
rect 196768 148102 197088 148170
rect 196768 148046 196838 148102
rect 196894 148046 196962 148102
rect 197018 148046 197088 148102
rect 196768 147978 197088 148046
rect 196768 147922 196838 147978
rect 196894 147922 196962 147978
rect 197018 147922 197088 147978
rect 196768 147888 197088 147922
rect 227488 148350 227808 148384
rect 227488 148294 227558 148350
rect 227614 148294 227682 148350
rect 227738 148294 227808 148350
rect 227488 148226 227808 148294
rect 227488 148170 227558 148226
rect 227614 148170 227682 148226
rect 227738 148170 227808 148226
rect 227488 148102 227808 148170
rect 227488 148046 227558 148102
rect 227614 148046 227682 148102
rect 227738 148046 227808 148102
rect 227488 147978 227808 148046
rect 227488 147922 227558 147978
rect 227614 147922 227682 147978
rect 227738 147922 227808 147978
rect 227488 147888 227808 147922
rect 258208 148350 258528 148384
rect 258208 148294 258278 148350
rect 258334 148294 258402 148350
rect 258458 148294 258528 148350
rect 258208 148226 258528 148294
rect 258208 148170 258278 148226
rect 258334 148170 258402 148226
rect 258458 148170 258528 148226
rect 258208 148102 258528 148170
rect 258208 148046 258278 148102
rect 258334 148046 258402 148102
rect 258458 148046 258528 148102
rect 258208 147978 258528 148046
rect 258208 147922 258278 147978
rect 258334 147922 258402 147978
rect 258458 147922 258528 147978
rect 258208 147888 258528 147922
rect 288928 148350 289248 148384
rect 288928 148294 288998 148350
rect 289054 148294 289122 148350
rect 289178 148294 289248 148350
rect 288928 148226 289248 148294
rect 288928 148170 288998 148226
rect 289054 148170 289122 148226
rect 289178 148170 289248 148226
rect 288928 148102 289248 148170
rect 288928 148046 288998 148102
rect 289054 148046 289122 148102
rect 289178 148046 289248 148102
rect 288928 147978 289248 148046
rect 288928 147922 288998 147978
rect 289054 147922 289122 147978
rect 289178 147922 289248 147978
rect 288928 147888 289248 147922
rect 319648 148350 319968 148384
rect 319648 148294 319718 148350
rect 319774 148294 319842 148350
rect 319898 148294 319968 148350
rect 319648 148226 319968 148294
rect 319648 148170 319718 148226
rect 319774 148170 319842 148226
rect 319898 148170 319968 148226
rect 319648 148102 319968 148170
rect 319648 148046 319718 148102
rect 319774 148046 319842 148102
rect 319898 148046 319968 148102
rect 319648 147978 319968 148046
rect 319648 147922 319718 147978
rect 319774 147922 319842 147978
rect 319898 147922 319968 147978
rect 319648 147888 319968 147922
rect 350368 148350 350688 148384
rect 350368 148294 350438 148350
rect 350494 148294 350562 148350
rect 350618 148294 350688 148350
rect 350368 148226 350688 148294
rect 350368 148170 350438 148226
rect 350494 148170 350562 148226
rect 350618 148170 350688 148226
rect 350368 148102 350688 148170
rect 350368 148046 350438 148102
rect 350494 148046 350562 148102
rect 350618 148046 350688 148102
rect 350368 147978 350688 148046
rect 350368 147922 350438 147978
rect 350494 147922 350562 147978
rect 350618 147922 350688 147978
rect 350368 147888 350688 147922
rect 381088 148350 381408 148384
rect 381088 148294 381158 148350
rect 381214 148294 381282 148350
rect 381338 148294 381408 148350
rect 381088 148226 381408 148294
rect 381088 148170 381158 148226
rect 381214 148170 381282 148226
rect 381338 148170 381408 148226
rect 381088 148102 381408 148170
rect 381088 148046 381158 148102
rect 381214 148046 381282 148102
rect 381338 148046 381408 148102
rect 381088 147978 381408 148046
rect 381088 147922 381158 147978
rect 381214 147922 381282 147978
rect 381338 147922 381408 147978
rect 381088 147888 381408 147922
rect 411808 148350 412128 148384
rect 411808 148294 411878 148350
rect 411934 148294 412002 148350
rect 412058 148294 412128 148350
rect 411808 148226 412128 148294
rect 411808 148170 411878 148226
rect 411934 148170 412002 148226
rect 412058 148170 412128 148226
rect 411808 148102 412128 148170
rect 411808 148046 411878 148102
rect 411934 148046 412002 148102
rect 412058 148046 412128 148102
rect 411808 147978 412128 148046
rect 411808 147922 411878 147978
rect 411934 147922 412002 147978
rect 412058 147922 412128 147978
rect 411808 147888 412128 147922
rect 442528 148350 442848 148384
rect 442528 148294 442598 148350
rect 442654 148294 442722 148350
rect 442778 148294 442848 148350
rect 442528 148226 442848 148294
rect 442528 148170 442598 148226
rect 442654 148170 442722 148226
rect 442778 148170 442848 148226
rect 442528 148102 442848 148170
rect 442528 148046 442598 148102
rect 442654 148046 442722 148102
rect 442778 148046 442848 148102
rect 442528 147978 442848 148046
rect 442528 147922 442598 147978
rect 442654 147922 442722 147978
rect 442778 147922 442848 147978
rect 442528 147888 442848 147922
rect 473248 148350 473568 148384
rect 473248 148294 473318 148350
rect 473374 148294 473442 148350
rect 473498 148294 473568 148350
rect 473248 148226 473568 148294
rect 473248 148170 473318 148226
rect 473374 148170 473442 148226
rect 473498 148170 473568 148226
rect 473248 148102 473568 148170
rect 473248 148046 473318 148102
rect 473374 148046 473442 148102
rect 473498 148046 473568 148102
rect 473248 147978 473568 148046
rect 473248 147922 473318 147978
rect 473374 147922 473442 147978
rect 473498 147922 473568 147978
rect 473248 147888 473568 147922
rect 503968 148350 504288 148384
rect 503968 148294 504038 148350
rect 504094 148294 504162 148350
rect 504218 148294 504288 148350
rect 503968 148226 504288 148294
rect 503968 148170 504038 148226
rect 504094 148170 504162 148226
rect 504218 148170 504288 148226
rect 503968 148102 504288 148170
rect 503968 148046 504038 148102
rect 504094 148046 504162 148102
rect 504218 148046 504288 148102
rect 503968 147978 504288 148046
rect 503968 147922 504038 147978
rect 504094 147922 504162 147978
rect 504218 147922 504288 147978
rect 503968 147888 504288 147922
rect 534688 148350 535008 148384
rect 534688 148294 534758 148350
rect 534814 148294 534882 148350
rect 534938 148294 535008 148350
rect 534688 148226 535008 148294
rect 534688 148170 534758 148226
rect 534814 148170 534882 148226
rect 534938 148170 535008 148226
rect 534688 148102 535008 148170
rect 534688 148046 534758 148102
rect 534814 148046 534882 148102
rect 534938 148046 535008 148102
rect 534688 147978 535008 148046
rect 534688 147922 534758 147978
rect 534814 147922 534882 147978
rect 534938 147922 535008 147978
rect 534688 147888 535008 147922
rect 565408 148350 565728 148384
rect 565408 148294 565478 148350
rect 565534 148294 565602 148350
rect 565658 148294 565728 148350
rect 565408 148226 565728 148294
rect 565408 148170 565478 148226
rect 565534 148170 565602 148226
rect 565658 148170 565728 148226
rect 565408 148102 565728 148170
rect 565408 148046 565478 148102
rect 565534 148046 565602 148102
rect 565658 148046 565728 148102
rect 565408 147978 565728 148046
rect 565408 147922 565478 147978
rect 565534 147922 565602 147978
rect 565658 147922 565728 147978
rect 565408 147888 565728 147922
rect 585452 146244 585508 165676
rect 585788 156996 585844 178892
rect 585788 156930 585844 156940
rect 589098 166350 589718 183922
rect 589098 166294 589194 166350
rect 589250 166294 589318 166350
rect 589374 166294 589442 166350
rect 589498 166294 589566 166350
rect 589622 166294 589718 166350
rect 589098 166226 589718 166294
rect 589098 166170 589194 166226
rect 589250 166170 589318 166226
rect 589374 166170 589442 166226
rect 589498 166170 589566 166226
rect 589622 166170 589718 166226
rect 589098 166102 589718 166170
rect 589098 166046 589194 166102
rect 589250 166046 589318 166102
rect 589374 166046 589442 166102
rect 589498 166046 589566 166102
rect 589622 166046 589718 166102
rect 589098 165978 589718 166046
rect 589098 165922 589194 165978
rect 589250 165922 589318 165978
rect 589374 165922 589442 165978
rect 589498 165922 589566 165978
rect 589622 165922 589718 165978
rect 585452 146178 585508 146188
rect 585564 152516 585620 152526
rect 6188 143938 6244 143948
rect 27808 136350 28128 136384
rect 27808 136294 27878 136350
rect 27934 136294 28002 136350
rect 28058 136294 28128 136350
rect 27808 136226 28128 136294
rect 27808 136170 27878 136226
rect 27934 136170 28002 136226
rect 28058 136170 28128 136226
rect 27808 136102 28128 136170
rect 27808 136046 27878 136102
rect 27934 136046 28002 136102
rect 28058 136046 28128 136102
rect 27808 135978 28128 136046
rect 27808 135922 27878 135978
rect 27934 135922 28002 135978
rect 28058 135922 28128 135978
rect 27808 135888 28128 135922
rect 58528 136350 58848 136384
rect 58528 136294 58598 136350
rect 58654 136294 58722 136350
rect 58778 136294 58848 136350
rect 58528 136226 58848 136294
rect 58528 136170 58598 136226
rect 58654 136170 58722 136226
rect 58778 136170 58848 136226
rect 58528 136102 58848 136170
rect 58528 136046 58598 136102
rect 58654 136046 58722 136102
rect 58778 136046 58848 136102
rect 58528 135978 58848 136046
rect 58528 135922 58598 135978
rect 58654 135922 58722 135978
rect 58778 135922 58848 135978
rect 58528 135888 58848 135922
rect 89248 136350 89568 136384
rect 89248 136294 89318 136350
rect 89374 136294 89442 136350
rect 89498 136294 89568 136350
rect 89248 136226 89568 136294
rect 89248 136170 89318 136226
rect 89374 136170 89442 136226
rect 89498 136170 89568 136226
rect 89248 136102 89568 136170
rect 89248 136046 89318 136102
rect 89374 136046 89442 136102
rect 89498 136046 89568 136102
rect 89248 135978 89568 136046
rect 89248 135922 89318 135978
rect 89374 135922 89442 135978
rect 89498 135922 89568 135978
rect 89248 135888 89568 135922
rect 119968 136350 120288 136384
rect 119968 136294 120038 136350
rect 120094 136294 120162 136350
rect 120218 136294 120288 136350
rect 119968 136226 120288 136294
rect 119968 136170 120038 136226
rect 120094 136170 120162 136226
rect 120218 136170 120288 136226
rect 119968 136102 120288 136170
rect 119968 136046 120038 136102
rect 120094 136046 120162 136102
rect 120218 136046 120288 136102
rect 119968 135978 120288 136046
rect 119968 135922 120038 135978
rect 120094 135922 120162 135978
rect 120218 135922 120288 135978
rect 119968 135888 120288 135922
rect 150688 136350 151008 136384
rect 150688 136294 150758 136350
rect 150814 136294 150882 136350
rect 150938 136294 151008 136350
rect 150688 136226 151008 136294
rect 150688 136170 150758 136226
rect 150814 136170 150882 136226
rect 150938 136170 151008 136226
rect 150688 136102 151008 136170
rect 150688 136046 150758 136102
rect 150814 136046 150882 136102
rect 150938 136046 151008 136102
rect 150688 135978 151008 136046
rect 150688 135922 150758 135978
rect 150814 135922 150882 135978
rect 150938 135922 151008 135978
rect 150688 135888 151008 135922
rect 181408 136350 181728 136384
rect 181408 136294 181478 136350
rect 181534 136294 181602 136350
rect 181658 136294 181728 136350
rect 181408 136226 181728 136294
rect 181408 136170 181478 136226
rect 181534 136170 181602 136226
rect 181658 136170 181728 136226
rect 181408 136102 181728 136170
rect 181408 136046 181478 136102
rect 181534 136046 181602 136102
rect 181658 136046 181728 136102
rect 181408 135978 181728 136046
rect 181408 135922 181478 135978
rect 181534 135922 181602 135978
rect 181658 135922 181728 135978
rect 181408 135888 181728 135922
rect 212128 136350 212448 136384
rect 212128 136294 212198 136350
rect 212254 136294 212322 136350
rect 212378 136294 212448 136350
rect 212128 136226 212448 136294
rect 212128 136170 212198 136226
rect 212254 136170 212322 136226
rect 212378 136170 212448 136226
rect 212128 136102 212448 136170
rect 212128 136046 212198 136102
rect 212254 136046 212322 136102
rect 212378 136046 212448 136102
rect 212128 135978 212448 136046
rect 212128 135922 212198 135978
rect 212254 135922 212322 135978
rect 212378 135922 212448 135978
rect 212128 135888 212448 135922
rect 242848 136350 243168 136384
rect 242848 136294 242918 136350
rect 242974 136294 243042 136350
rect 243098 136294 243168 136350
rect 242848 136226 243168 136294
rect 242848 136170 242918 136226
rect 242974 136170 243042 136226
rect 243098 136170 243168 136226
rect 242848 136102 243168 136170
rect 242848 136046 242918 136102
rect 242974 136046 243042 136102
rect 243098 136046 243168 136102
rect 242848 135978 243168 136046
rect 242848 135922 242918 135978
rect 242974 135922 243042 135978
rect 243098 135922 243168 135978
rect 242848 135888 243168 135922
rect 273568 136350 273888 136384
rect 273568 136294 273638 136350
rect 273694 136294 273762 136350
rect 273818 136294 273888 136350
rect 273568 136226 273888 136294
rect 273568 136170 273638 136226
rect 273694 136170 273762 136226
rect 273818 136170 273888 136226
rect 273568 136102 273888 136170
rect 273568 136046 273638 136102
rect 273694 136046 273762 136102
rect 273818 136046 273888 136102
rect 273568 135978 273888 136046
rect 273568 135922 273638 135978
rect 273694 135922 273762 135978
rect 273818 135922 273888 135978
rect 273568 135888 273888 135922
rect 304288 136350 304608 136384
rect 304288 136294 304358 136350
rect 304414 136294 304482 136350
rect 304538 136294 304608 136350
rect 304288 136226 304608 136294
rect 304288 136170 304358 136226
rect 304414 136170 304482 136226
rect 304538 136170 304608 136226
rect 304288 136102 304608 136170
rect 304288 136046 304358 136102
rect 304414 136046 304482 136102
rect 304538 136046 304608 136102
rect 304288 135978 304608 136046
rect 304288 135922 304358 135978
rect 304414 135922 304482 135978
rect 304538 135922 304608 135978
rect 304288 135888 304608 135922
rect 335008 136350 335328 136384
rect 335008 136294 335078 136350
rect 335134 136294 335202 136350
rect 335258 136294 335328 136350
rect 335008 136226 335328 136294
rect 335008 136170 335078 136226
rect 335134 136170 335202 136226
rect 335258 136170 335328 136226
rect 335008 136102 335328 136170
rect 335008 136046 335078 136102
rect 335134 136046 335202 136102
rect 335258 136046 335328 136102
rect 335008 135978 335328 136046
rect 335008 135922 335078 135978
rect 335134 135922 335202 135978
rect 335258 135922 335328 135978
rect 335008 135888 335328 135922
rect 365728 136350 366048 136384
rect 365728 136294 365798 136350
rect 365854 136294 365922 136350
rect 365978 136294 366048 136350
rect 365728 136226 366048 136294
rect 365728 136170 365798 136226
rect 365854 136170 365922 136226
rect 365978 136170 366048 136226
rect 365728 136102 366048 136170
rect 365728 136046 365798 136102
rect 365854 136046 365922 136102
rect 365978 136046 366048 136102
rect 365728 135978 366048 136046
rect 365728 135922 365798 135978
rect 365854 135922 365922 135978
rect 365978 135922 366048 135978
rect 365728 135888 366048 135922
rect 396448 136350 396768 136384
rect 396448 136294 396518 136350
rect 396574 136294 396642 136350
rect 396698 136294 396768 136350
rect 396448 136226 396768 136294
rect 396448 136170 396518 136226
rect 396574 136170 396642 136226
rect 396698 136170 396768 136226
rect 396448 136102 396768 136170
rect 396448 136046 396518 136102
rect 396574 136046 396642 136102
rect 396698 136046 396768 136102
rect 396448 135978 396768 136046
rect 396448 135922 396518 135978
rect 396574 135922 396642 135978
rect 396698 135922 396768 135978
rect 396448 135888 396768 135922
rect 427168 136350 427488 136384
rect 427168 136294 427238 136350
rect 427294 136294 427362 136350
rect 427418 136294 427488 136350
rect 427168 136226 427488 136294
rect 427168 136170 427238 136226
rect 427294 136170 427362 136226
rect 427418 136170 427488 136226
rect 427168 136102 427488 136170
rect 427168 136046 427238 136102
rect 427294 136046 427362 136102
rect 427418 136046 427488 136102
rect 427168 135978 427488 136046
rect 427168 135922 427238 135978
rect 427294 135922 427362 135978
rect 427418 135922 427488 135978
rect 427168 135888 427488 135922
rect 457888 136350 458208 136384
rect 457888 136294 457958 136350
rect 458014 136294 458082 136350
rect 458138 136294 458208 136350
rect 457888 136226 458208 136294
rect 457888 136170 457958 136226
rect 458014 136170 458082 136226
rect 458138 136170 458208 136226
rect 457888 136102 458208 136170
rect 457888 136046 457958 136102
rect 458014 136046 458082 136102
rect 458138 136046 458208 136102
rect 457888 135978 458208 136046
rect 457888 135922 457958 135978
rect 458014 135922 458082 135978
rect 458138 135922 458208 135978
rect 457888 135888 458208 135922
rect 488608 136350 488928 136384
rect 488608 136294 488678 136350
rect 488734 136294 488802 136350
rect 488858 136294 488928 136350
rect 488608 136226 488928 136294
rect 488608 136170 488678 136226
rect 488734 136170 488802 136226
rect 488858 136170 488928 136226
rect 488608 136102 488928 136170
rect 488608 136046 488678 136102
rect 488734 136046 488802 136102
rect 488858 136046 488928 136102
rect 488608 135978 488928 136046
rect 488608 135922 488678 135978
rect 488734 135922 488802 135978
rect 488858 135922 488928 135978
rect 488608 135888 488928 135922
rect 519328 136350 519648 136384
rect 519328 136294 519398 136350
rect 519454 136294 519522 136350
rect 519578 136294 519648 136350
rect 519328 136226 519648 136294
rect 519328 136170 519398 136226
rect 519454 136170 519522 136226
rect 519578 136170 519648 136226
rect 519328 136102 519648 136170
rect 519328 136046 519398 136102
rect 519454 136046 519522 136102
rect 519578 136046 519648 136102
rect 519328 135978 519648 136046
rect 519328 135922 519398 135978
rect 519454 135922 519522 135978
rect 519578 135922 519648 135978
rect 519328 135888 519648 135922
rect 550048 136350 550368 136384
rect 550048 136294 550118 136350
rect 550174 136294 550242 136350
rect 550298 136294 550368 136350
rect 550048 136226 550368 136294
rect 550048 136170 550118 136226
rect 550174 136170 550242 136226
rect 550298 136170 550368 136226
rect 550048 136102 550368 136170
rect 550048 136046 550118 136102
rect 550174 136046 550242 136102
rect 550298 136046 550368 136102
rect 550048 135978 550368 136046
rect 550048 135922 550118 135978
rect 550174 135922 550242 135978
rect 550298 135922 550368 135978
rect 550048 135888 550368 135922
rect 585564 135492 585620 152460
rect 585564 135426 585620 135436
rect 589098 148350 589718 165922
rect 589098 148294 589194 148350
rect 589250 148294 589318 148350
rect 589374 148294 589442 148350
rect 589498 148294 589566 148350
rect 589622 148294 589718 148350
rect 589098 148226 589718 148294
rect 589098 148170 589194 148226
rect 589250 148170 589318 148226
rect 589374 148170 589442 148226
rect 589498 148170 589566 148226
rect 589622 148170 589718 148226
rect 589098 148102 589718 148170
rect 589098 148046 589194 148102
rect 589250 148046 589318 148102
rect 589374 148046 589442 148102
rect 589498 148046 589566 148102
rect 589622 148046 589718 148102
rect 589098 147978 589718 148046
rect 589098 147922 589194 147978
rect 589250 147922 589318 147978
rect 589374 147922 589442 147978
rect 589498 147922 589566 147978
rect 589622 147922 589718 147978
rect 5418 130294 5514 130350
rect 5570 130294 5638 130350
rect 5694 130294 5762 130350
rect 5818 130294 5886 130350
rect 5942 130294 6038 130350
rect 5418 130226 6038 130294
rect 5418 130170 5514 130226
rect 5570 130170 5638 130226
rect 5694 130170 5762 130226
rect 5818 130170 5886 130226
rect 5942 130170 6038 130226
rect 5418 130102 6038 130170
rect 5418 130046 5514 130102
rect 5570 130046 5638 130102
rect 5694 130046 5762 130102
rect 5818 130046 5886 130102
rect 5942 130046 6038 130102
rect 5418 129978 6038 130046
rect 5418 129922 5514 129978
rect 5570 129922 5638 129978
rect 5694 129922 5762 129978
rect 5818 129922 5886 129978
rect 5942 129922 6038 129978
rect -956 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 -336 112350
rect -956 112226 -336 112294
rect -956 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 -336 112226
rect -956 112102 -336 112170
rect -956 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 -336 112102
rect -956 111978 -336 112046
rect -956 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 -336 111978
rect -956 94350 -336 111922
rect 4172 121492 4228 121502
rect 4172 101892 4228 121436
rect 4172 101826 4228 101836
rect 5418 112350 6038 129922
rect 12448 130350 12768 130384
rect 12448 130294 12518 130350
rect 12574 130294 12642 130350
rect 12698 130294 12768 130350
rect 12448 130226 12768 130294
rect 12448 130170 12518 130226
rect 12574 130170 12642 130226
rect 12698 130170 12768 130226
rect 12448 130102 12768 130170
rect 12448 130046 12518 130102
rect 12574 130046 12642 130102
rect 12698 130046 12768 130102
rect 12448 129978 12768 130046
rect 12448 129922 12518 129978
rect 12574 129922 12642 129978
rect 12698 129922 12768 129978
rect 12448 129888 12768 129922
rect 43168 130350 43488 130384
rect 43168 130294 43238 130350
rect 43294 130294 43362 130350
rect 43418 130294 43488 130350
rect 43168 130226 43488 130294
rect 43168 130170 43238 130226
rect 43294 130170 43362 130226
rect 43418 130170 43488 130226
rect 43168 130102 43488 130170
rect 43168 130046 43238 130102
rect 43294 130046 43362 130102
rect 43418 130046 43488 130102
rect 43168 129978 43488 130046
rect 43168 129922 43238 129978
rect 43294 129922 43362 129978
rect 43418 129922 43488 129978
rect 43168 129888 43488 129922
rect 73888 130350 74208 130384
rect 73888 130294 73958 130350
rect 74014 130294 74082 130350
rect 74138 130294 74208 130350
rect 73888 130226 74208 130294
rect 73888 130170 73958 130226
rect 74014 130170 74082 130226
rect 74138 130170 74208 130226
rect 73888 130102 74208 130170
rect 73888 130046 73958 130102
rect 74014 130046 74082 130102
rect 74138 130046 74208 130102
rect 73888 129978 74208 130046
rect 73888 129922 73958 129978
rect 74014 129922 74082 129978
rect 74138 129922 74208 129978
rect 73888 129888 74208 129922
rect 104608 130350 104928 130384
rect 104608 130294 104678 130350
rect 104734 130294 104802 130350
rect 104858 130294 104928 130350
rect 104608 130226 104928 130294
rect 104608 130170 104678 130226
rect 104734 130170 104802 130226
rect 104858 130170 104928 130226
rect 104608 130102 104928 130170
rect 104608 130046 104678 130102
rect 104734 130046 104802 130102
rect 104858 130046 104928 130102
rect 104608 129978 104928 130046
rect 104608 129922 104678 129978
rect 104734 129922 104802 129978
rect 104858 129922 104928 129978
rect 104608 129888 104928 129922
rect 135328 130350 135648 130384
rect 135328 130294 135398 130350
rect 135454 130294 135522 130350
rect 135578 130294 135648 130350
rect 135328 130226 135648 130294
rect 135328 130170 135398 130226
rect 135454 130170 135522 130226
rect 135578 130170 135648 130226
rect 135328 130102 135648 130170
rect 135328 130046 135398 130102
rect 135454 130046 135522 130102
rect 135578 130046 135648 130102
rect 135328 129978 135648 130046
rect 135328 129922 135398 129978
rect 135454 129922 135522 129978
rect 135578 129922 135648 129978
rect 135328 129888 135648 129922
rect 166048 130350 166368 130384
rect 166048 130294 166118 130350
rect 166174 130294 166242 130350
rect 166298 130294 166368 130350
rect 166048 130226 166368 130294
rect 166048 130170 166118 130226
rect 166174 130170 166242 130226
rect 166298 130170 166368 130226
rect 166048 130102 166368 130170
rect 166048 130046 166118 130102
rect 166174 130046 166242 130102
rect 166298 130046 166368 130102
rect 166048 129978 166368 130046
rect 166048 129922 166118 129978
rect 166174 129922 166242 129978
rect 166298 129922 166368 129978
rect 166048 129888 166368 129922
rect 196768 130350 197088 130384
rect 196768 130294 196838 130350
rect 196894 130294 196962 130350
rect 197018 130294 197088 130350
rect 196768 130226 197088 130294
rect 196768 130170 196838 130226
rect 196894 130170 196962 130226
rect 197018 130170 197088 130226
rect 196768 130102 197088 130170
rect 196768 130046 196838 130102
rect 196894 130046 196962 130102
rect 197018 130046 197088 130102
rect 196768 129978 197088 130046
rect 196768 129922 196838 129978
rect 196894 129922 196962 129978
rect 197018 129922 197088 129978
rect 196768 129888 197088 129922
rect 227488 130350 227808 130384
rect 227488 130294 227558 130350
rect 227614 130294 227682 130350
rect 227738 130294 227808 130350
rect 227488 130226 227808 130294
rect 227488 130170 227558 130226
rect 227614 130170 227682 130226
rect 227738 130170 227808 130226
rect 227488 130102 227808 130170
rect 227488 130046 227558 130102
rect 227614 130046 227682 130102
rect 227738 130046 227808 130102
rect 227488 129978 227808 130046
rect 227488 129922 227558 129978
rect 227614 129922 227682 129978
rect 227738 129922 227808 129978
rect 227488 129888 227808 129922
rect 258208 130350 258528 130384
rect 258208 130294 258278 130350
rect 258334 130294 258402 130350
rect 258458 130294 258528 130350
rect 258208 130226 258528 130294
rect 258208 130170 258278 130226
rect 258334 130170 258402 130226
rect 258458 130170 258528 130226
rect 258208 130102 258528 130170
rect 258208 130046 258278 130102
rect 258334 130046 258402 130102
rect 258458 130046 258528 130102
rect 258208 129978 258528 130046
rect 258208 129922 258278 129978
rect 258334 129922 258402 129978
rect 258458 129922 258528 129978
rect 258208 129888 258528 129922
rect 288928 130350 289248 130384
rect 288928 130294 288998 130350
rect 289054 130294 289122 130350
rect 289178 130294 289248 130350
rect 288928 130226 289248 130294
rect 288928 130170 288998 130226
rect 289054 130170 289122 130226
rect 289178 130170 289248 130226
rect 288928 130102 289248 130170
rect 288928 130046 288998 130102
rect 289054 130046 289122 130102
rect 289178 130046 289248 130102
rect 288928 129978 289248 130046
rect 288928 129922 288998 129978
rect 289054 129922 289122 129978
rect 289178 129922 289248 129978
rect 288928 129888 289248 129922
rect 319648 130350 319968 130384
rect 319648 130294 319718 130350
rect 319774 130294 319842 130350
rect 319898 130294 319968 130350
rect 319648 130226 319968 130294
rect 319648 130170 319718 130226
rect 319774 130170 319842 130226
rect 319898 130170 319968 130226
rect 319648 130102 319968 130170
rect 319648 130046 319718 130102
rect 319774 130046 319842 130102
rect 319898 130046 319968 130102
rect 319648 129978 319968 130046
rect 319648 129922 319718 129978
rect 319774 129922 319842 129978
rect 319898 129922 319968 129978
rect 319648 129888 319968 129922
rect 350368 130350 350688 130384
rect 350368 130294 350438 130350
rect 350494 130294 350562 130350
rect 350618 130294 350688 130350
rect 350368 130226 350688 130294
rect 350368 130170 350438 130226
rect 350494 130170 350562 130226
rect 350618 130170 350688 130226
rect 350368 130102 350688 130170
rect 350368 130046 350438 130102
rect 350494 130046 350562 130102
rect 350618 130046 350688 130102
rect 350368 129978 350688 130046
rect 350368 129922 350438 129978
rect 350494 129922 350562 129978
rect 350618 129922 350688 129978
rect 350368 129888 350688 129922
rect 381088 130350 381408 130384
rect 381088 130294 381158 130350
rect 381214 130294 381282 130350
rect 381338 130294 381408 130350
rect 381088 130226 381408 130294
rect 381088 130170 381158 130226
rect 381214 130170 381282 130226
rect 381338 130170 381408 130226
rect 381088 130102 381408 130170
rect 381088 130046 381158 130102
rect 381214 130046 381282 130102
rect 381338 130046 381408 130102
rect 381088 129978 381408 130046
rect 381088 129922 381158 129978
rect 381214 129922 381282 129978
rect 381338 129922 381408 129978
rect 381088 129888 381408 129922
rect 411808 130350 412128 130384
rect 411808 130294 411878 130350
rect 411934 130294 412002 130350
rect 412058 130294 412128 130350
rect 411808 130226 412128 130294
rect 411808 130170 411878 130226
rect 411934 130170 412002 130226
rect 412058 130170 412128 130226
rect 411808 130102 412128 130170
rect 411808 130046 411878 130102
rect 411934 130046 412002 130102
rect 412058 130046 412128 130102
rect 411808 129978 412128 130046
rect 411808 129922 411878 129978
rect 411934 129922 412002 129978
rect 412058 129922 412128 129978
rect 411808 129888 412128 129922
rect 442528 130350 442848 130384
rect 442528 130294 442598 130350
rect 442654 130294 442722 130350
rect 442778 130294 442848 130350
rect 442528 130226 442848 130294
rect 442528 130170 442598 130226
rect 442654 130170 442722 130226
rect 442778 130170 442848 130226
rect 442528 130102 442848 130170
rect 442528 130046 442598 130102
rect 442654 130046 442722 130102
rect 442778 130046 442848 130102
rect 442528 129978 442848 130046
rect 442528 129922 442598 129978
rect 442654 129922 442722 129978
rect 442778 129922 442848 129978
rect 442528 129888 442848 129922
rect 473248 130350 473568 130384
rect 473248 130294 473318 130350
rect 473374 130294 473442 130350
rect 473498 130294 473568 130350
rect 473248 130226 473568 130294
rect 473248 130170 473318 130226
rect 473374 130170 473442 130226
rect 473498 130170 473568 130226
rect 473248 130102 473568 130170
rect 473248 130046 473318 130102
rect 473374 130046 473442 130102
rect 473498 130046 473568 130102
rect 473248 129978 473568 130046
rect 473248 129922 473318 129978
rect 473374 129922 473442 129978
rect 473498 129922 473568 129978
rect 473248 129888 473568 129922
rect 503968 130350 504288 130384
rect 503968 130294 504038 130350
rect 504094 130294 504162 130350
rect 504218 130294 504288 130350
rect 503968 130226 504288 130294
rect 503968 130170 504038 130226
rect 504094 130170 504162 130226
rect 504218 130170 504288 130226
rect 503968 130102 504288 130170
rect 503968 130046 504038 130102
rect 504094 130046 504162 130102
rect 504218 130046 504288 130102
rect 503968 129978 504288 130046
rect 503968 129922 504038 129978
rect 504094 129922 504162 129978
rect 504218 129922 504288 129978
rect 503968 129888 504288 129922
rect 534688 130350 535008 130384
rect 534688 130294 534758 130350
rect 534814 130294 534882 130350
rect 534938 130294 535008 130350
rect 534688 130226 535008 130294
rect 534688 130170 534758 130226
rect 534814 130170 534882 130226
rect 534938 130170 535008 130226
rect 534688 130102 535008 130170
rect 534688 130046 534758 130102
rect 534814 130046 534882 130102
rect 534938 130046 535008 130102
rect 534688 129978 535008 130046
rect 534688 129922 534758 129978
rect 534814 129922 534882 129978
rect 534938 129922 535008 129978
rect 534688 129888 535008 129922
rect 565408 130350 565728 130384
rect 565408 130294 565478 130350
rect 565534 130294 565602 130350
rect 565658 130294 565728 130350
rect 565408 130226 565728 130294
rect 565408 130170 565478 130226
rect 565534 130170 565602 130226
rect 565658 130170 565728 130226
rect 565408 130102 565728 130170
rect 565408 130046 565478 130102
rect 565534 130046 565602 130102
rect 565658 130046 565728 130102
rect 565408 129978 565728 130046
rect 565408 129922 565478 129978
rect 565534 129922 565602 129978
rect 565658 129922 565728 129978
rect 565408 129888 565728 129922
rect 589098 130350 589718 147922
rect 592818 208350 593438 225922
rect 592818 208294 592914 208350
rect 592970 208294 593038 208350
rect 593094 208294 593162 208350
rect 593218 208294 593286 208350
rect 593342 208294 593438 208350
rect 592818 208226 593438 208294
rect 592818 208170 592914 208226
rect 592970 208170 593038 208226
rect 593094 208170 593162 208226
rect 593218 208170 593286 208226
rect 593342 208170 593438 208226
rect 592818 208102 593438 208170
rect 592818 208046 592914 208102
rect 592970 208046 593038 208102
rect 593094 208046 593162 208102
rect 593218 208046 593286 208102
rect 593342 208046 593438 208102
rect 592818 207978 593438 208046
rect 592818 207922 592914 207978
rect 592970 207922 593038 207978
rect 593094 207922 593162 207978
rect 593218 207922 593286 207978
rect 593342 207922 593438 207978
rect 592818 190350 593438 207922
rect 592818 190294 592914 190350
rect 592970 190294 593038 190350
rect 593094 190294 593162 190350
rect 593218 190294 593286 190350
rect 593342 190294 593438 190350
rect 592818 190226 593438 190294
rect 592818 190170 592914 190226
rect 592970 190170 593038 190226
rect 593094 190170 593162 190226
rect 593218 190170 593286 190226
rect 593342 190170 593438 190226
rect 592818 190102 593438 190170
rect 592818 190046 592914 190102
rect 592970 190046 593038 190102
rect 593094 190046 593162 190102
rect 593218 190046 593286 190102
rect 593342 190046 593438 190102
rect 592818 189978 593438 190046
rect 592818 189922 592914 189978
rect 592970 189922 593038 189978
rect 593094 189922 593162 189978
rect 593218 189922 593286 189978
rect 593342 189922 593438 189978
rect 592818 172350 593438 189922
rect 592818 172294 592914 172350
rect 592970 172294 593038 172350
rect 593094 172294 593162 172350
rect 593218 172294 593286 172350
rect 593342 172294 593438 172350
rect 592818 172226 593438 172294
rect 592818 172170 592914 172226
rect 592970 172170 593038 172226
rect 593094 172170 593162 172226
rect 593218 172170 593286 172226
rect 593342 172170 593438 172226
rect 592818 172102 593438 172170
rect 592818 172046 592914 172102
rect 592970 172046 593038 172102
rect 593094 172046 593162 172102
rect 593218 172046 593286 172102
rect 593342 172046 593438 172102
rect 592818 171978 593438 172046
rect 592818 171922 592914 171978
rect 592970 171922 593038 171978
rect 593094 171922 593162 171978
rect 593218 171922 593286 171978
rect 593342 171922 593438 171978
rect 592818 154350 593438 171922
rect 592818 154294 592914 154350
rect 592970 154294 593038 154350
rect 593094 154294 593162 154350
rect 593218 154294 593286 154350
rect 593342 154294 593438 154350
rect 592818 154226 593438 154294
rect 592818 154170 592914 154226
rect 592970 154170 593038 154226
rect 593094 154170 593162 154226
rect 593218 154170 593286 154226
rect 593342 154170 593438 154226
rect 592818 154102 593438 154170
rect 592818 154046 592914 154102
rect 592970 154046 593038 154102
rect 593094 154046 593162 154102
rect 593218 154046 593286 154102
rect 593342 154046 593438 154102
rect 592818 153978 593438 154046
rect 592818 153922 592914 153978
rect 592970 153922 593038 153978
rect 593094 153922 593162 153978
rect 593218 153922 593286 153978
rect 593342 153922 593438 153978
rect 589098 130294 589194 130350
rect 589250 130294 589318 130350
rect 589374 130294 589442 130350
rect 589498 130294 589566 130350
rect 589622 130294 589718 130350
rect 589098 130226 589718 130294
rect 589098 130170 589194 130226
rect 589250 130170 589318 130226
rect 589374 130170 589442 130226
rect 589498 130170 589566 130226
rect 589622 130170 589718 130226
rect 589098 130102 589718 130170
rect 589098 130046 589194 130102
rect 589250 130046 589318 130102
rect 589374 130046 589442 130102
rect 589498 130046 589566 130102
rect 589622 130046 589718 130102
rect 589098 129978 589718 130046
rect 589098 129922 589194 129978
rect 589250 129922 589318 129978
rect 589374 129922 589442 129978
rect 589498 129922 589566 129978
rect 589622 129922 589718 129978
rect 27808 118350 28128 118384
rect 27808 118294 27878 118350
rect 27934 118294 28002 118350
rect 28058 118294 28128 118350
rect 27808 118226 28128 118294
rect 27808 118170 27878 118226
rect 27934 118170 28002 118226
rect 28058 118170 28128 118226
rect 27808 118102 28128 118170
rect 27808 118046 27878 118102
rect 27934 118046 28002 118102
rect 28058 118046 28128 118102
rect 27808 117978 28128 118046
rect 27808 117922 27878 117978
rect 27934 117922 28002 117978
rect 28058 117922 28128 117978
rect 27808 117888 28128 117922
rect 58528 118350 58848 118384
rect 58528 118294 58598 118350
rect 58654 118294 58722 118350
rect 58778 118294 58848 118350
rect 58528 118226 58848 118294
rect 58528 118170 58598 118226
rect 58654 118170 58722 118226
rect 58778 118170 58848 118226
rect 58528 118102 58848 118170
rect 58528 118046 58598 118102
rect 58654 118046 58722 118102
rect 58778 118046 58848 118102
rect 58528 117978 58848 118046
rect 58528 117922 58598 117978
rect 58654 117922 58722 117978
rect 58778 117922 58848 117978
rect 58528 117888 58848 117922
rect 89248 118350 89568 118384
rect 89248 118294 89318 118350
rect 89374 118294 89442 118350
rect 89498 118294 89568 118350
rect 89248 118226 89568 118294
rect 89248 118170 89318 118226
rect 89374 118170 89442 118226
rect 89498 118170 89568 118226
rect 89248 118102 89568 118170
rect 89248 118046 89318 118102
rect 89374 118046 89442 118102
rect 89498 118046 89568 118102
rect 89248 117978 89568 118046
rect 89248 117922 89318 117978
rect 89374 117922 89442 117978
rect 89498 117922 89568 117978
rect 89248 117888 89568 117922
rect 119968 118350 120288 118384
rect 119968 118294 120038 118350
rect 120094 118294 120162 118350
rect 120218 118294 120288 118350
rect 119968 118226 120288 118294
rect 119968 118170 120038 118226
rect 120094 118170 120162 118226
rect 120218 118170 120288 118226
rect 119968 118102 120288 118170
rect 119968 118046 120038 118102
rect 120094 118046 120162 118102
rect 120218 118046 120288 118102
rect 119968 117978 120288 118046
rect 119968 117922 120038 117978
rect 120094 117922 120162 117978
rect 120218 117922 120288 117978
rect 119968 117888 120288 117922
rect 150688 118350 151008 118384
rect 150688 118294 150758 118350
rect 150814 118294 150882 118350
rect 150938 118294 151008 118350
rect 150688 118226 151008 118294
rect 150688 118170 150758 118226
rect 150814 118170 150882 118226
rect 150938 118170 151008 118226
rect 150688 118102 151008 118170
rect 150688 118046 150758 118102
rect 150814 118046 150882 118102
rect 150938 118046 151008 118102
rect 150688 117978 151008 118046
rect 150688 117922 150758 117978
rect 150814 117922 150882 117978
rect 150938 117922 151008 117978
rect 150688 117888 151008 117922
rect 181408 118350 181728 118384
rect 181408 118294 181478 118350
rect 181534 118294 181602 118350
rect 181658 118294 181728 118350
rect 181408 118226 181728 118294
rect 181408 118170 181478 118226
rect 181534 118170 181602 118226
rect 181658 118170 181728 118226
rect 181408 118102 181728 118170
rect 181408 118046 181478 118102
rect 181534 118046 181602 118102
rect 181658 118046 181728 118102
rect 181408 117978 181728 118046
rect 181408 117922 181478 117978
rect 181534 117922 181602 117978
rect 181658 117922 181728 117978
rect 181408 117888 181728 117922
rect 212128 118350 212448 118384
rect 212128 118294 212198 118350
rect 212254 118294 212322 118350
rect 212378 118294 212448 118350
rect 212128 118226 212448 118294
rect 212128 118170 212198 118226
rect 212254 118170 212322 118226
rect 212378 118170 212448 118226
rect 212128 118102 212448 118170
rect 212128 118046 212198 118102
rect 212254 118046 212322 118102
rect 212378 118046 212448 118102
rect 212128 117978 212448 118046
rect 212128 117922 212198 117978
rect 212254 117922 212322 117978
rect 212378 117922 212448 117978
rect 212128 117888 212448 117922
rect 242848 118350 243168 118384
rect 242848 118294 242918 118350
rect 242974 118294 243042 118350
rect 243098 118294 243168 118350
rect 242848 118226 243168 118294
rect 242848 118170 242918 118226
rect 242974 118170 243042 118226
rect 243098 118170 243168 118226
rect 242848 118102 243168 118170
rect 242848 118046 242918 118102
rect 242974 118046 243042 118102
rect 243098 118046 243168 118102
rect 242848 117978 243168 118046
rect 242848 117922 242918 117978
rect 242974 117922 243042 117978
rect 243098 117922 243168 117978
rect 242848 117888 243168 117922
rect 273568 118350 273888 118384
rect 273568 118294 273638 118350
rect 273694 118294 273762 118350
rect 273818 118294 273888 118350
rect 273568 118226 273888 118294
rect 273568 118170 273638 118226
rect 273694 118170 273762 118226
rect 273818 118170 273888 118226
rect 273568 118102 273888 118170
rect 273568 118046 273638 118102
rect 273694 118046 273762 118102
rect 273818 118046 273888 118102
rect 273568 117978 273888 118046
rect 273568 117922 273638 117978
rect 273694 117922 273762 117978
rect 273818 117922 273888 117978
rect 273568 117888 273888 117922
rect 304288 118350 304608 118384
rect 304288 118294 304358 118350
rect 304414 118294 304482 118350
rect 304538 118294 304608 118350
rect 304288 118226 304608 118294
rect 304288 118170 304358 118226
rect 304414 118170 304482 118226
rect 304538 118170 304608 118226
rect 304288 118102 304608 118170
rect 304288 118046 304358 118102
rect 304414 118046 304482 118102
rect 304538 118046 304608 118102
rect 304288 117978 304608 118046
rect 304288 117922 304358 117978
rect 304414 117922 304482 117978
rect 304538 117922 304608 117978
rect 304288 117888 304608 117922
rect 335008 118350 335328 118384
rect 335008 118294 335078 118350
rect 335134 118294 335202 118350
rect 335258 118294 335328 118350
rect 335008 118226 335328 118294
rect 335008 118170 335078 118226
rect 335134 118170 335202 118226
rect 335258 118170 335328 118226
rect 335008 118102 335328 118170
rect 335008 118046 335078 118102
rect 335134 118046 335202 118102
rect 335258 118046 335328 118102
rect 335008 117978 335328 118046
rect 335008 117922 335078 117978
rect 335134 117922 335202 117978
rect 335258 117922 335328 117978
rect 335008 117888 335328 117922
rect 365728 118350 366048 118384
rect 365728 118294 365798 118350
rect 365854 118294 365922 118350
rect 365978 118294 366048 118350
rect 365728 118226 366048 118294
rect 365728 118170 365798 118226
rect 365854 118170 365922 118226
rect 365978 118170 366048 118226
rect 365728 118102 366048 118170
rect 365728 118046 365798 118102
rect 365854 118046 365922 118102
rect 365978 118046 366048 118102
rect 365728 117978 366048 118046
rect 365728 117922 365798 117978
rect 365854 117922 365922 117978
rect 365978 117922 366048 117978
rect 365728 117888 366048 117922
rect 396448 118350 396768 118384
rect 396448 118294 396518 118350
rect 396574 118294 396642 118350
rect 396698 118294 396768 118350
rect 396448 118226 396768 118294
rect 396448 118170 396518 118226
rect 396574 118170 396642 118226
rect 396698 118170 396768 118226
rect 396448 118102 396768 118170
rect 396448 118046 396518 118102
rect 396574 118046 396642 118102
rect 396698 118046 396768 118102
rect 396448 117978 396768 118046
rect 396448 117922 396518 117978
rect 396574 117922 396642 117978
rect 396698 117922 396768 117978
rect 396448 117888 396768 117922
rect 427168 118350 427488 118384
rect 427168 118294 427238 118350
rect 427294 118294 427362 118350
rect 427418 118294 427488 118350
rect 427168 118226 427488 118294
rect 427168 118170 427238 118226
rect 427294 118170 427362 118226
rect 427418 118170 427488 118226
rect 427168 118102 427488 118170
rect 427168 118046 427238 118102
rect 427294 118046 427362 118102
rect 427418 118046 427488 118102
rect 427168 117978 427488 118046
rect 427168 117922 427238 117978
rect 427294 117922 427362 117978
rect 427418 117922 427488 117978
rect 427168 117888 427488 117922
rect 457888 118350 458208 118384
rect 457888 118294 457958 118350
rect 458014 118294 458082 118350
rect 458138 118294 458208 118350
rect 457888 118226 458208 118294
rect 457888 118170 457958 118226
rect 458014 118170 458082 118226
rect 458138 118170 458208 118226
rect 457888 118102 458208 118170
rect 457888 118046 457958 118102
rect 458014 118046 458082 118102
rect 458138 118046 458208 118102
rect 457888 117978 458208 118046
rect 457888 117922 457958 117978
rect 458014 117922 458082 117978
rect 458138 117922 458208 117978
rect 457888 117888 458208 117922
rect 488608 118350 488928 118384
rect 488608 118294 488678 118350
rect 488734 118294 488802 118350
rect 488858 118294 488928 118350
rect 488608 118226 488928 118294
rect 488608 118170 488678 118226
rect 488734 118170 488802 118226
rect 488858 118170 488928 118226
rect 488608 118102 488928 118170
rect 488608 118046 488678 118102
rect 488734 118046 488802 118102
rect 488858 118046 488928 118102
rect 488608 117978 488928 118046
rect 488608 117922 488678 117978
rect 488734 117922 488802 117978
rect 488858 117922 488928 117978
rect 488608 117888 488928 117922
rect 519328 118350 519648 118384
rect 519328 118294 519398 118350
rect 519454 118294 519522 118350
rect 519578 118294 519648 118350
rect 519328 118226 519648 118294
rect 519328 118170 519398 118226
rect 519454 118170 519522 118226
rect 519578 118170 519648 118226
rect 519328 118102 519648 118170
rect 519328 118046 519398 118102
rect 519454 118046 519522 118102
rect 519578 118046 519648 118102
rect 519328 117978 519648 118046
rect 519328 117922 519398 117978
rect 519454 117922 519522 117978
rect 519578 117922 519648 117978
rect 519328 117888 519648 117922
rect 550048 118350 550368 118384
rect 550048 118294 550118 118350
rect 550174 118294 550242 118350
rect 550298 118294 550368 118350
rect 550048 118226 550368 118294
rect 550048 118170 550118 118226
rect 550174 118170 550242 118226
rect 550298 118170 550368 118226
rect 550048 118102 550368 118170
rect 550048 118046 550118 118102
rect 550174 118046 550242 118102
rect 550298 118046 550368 118102
rect 550048 117978 550368 118046
rect 550048 117922 550118 117978
rect 550174 117922 550242 117978
rect 550298 117922 550368 117978
rect 550048 117888 550368 117922
rect 5418 112294 5514 112350
rect 5570 112294 5638 112350
rect 5694 112294 5762 112350
rect 5818 112294 5886 112350
rect 5942 112294 6038 112350
rect 5418 112226 6038 112294
rect 5418 112170 5514 112226
rect 5570 112170 5638 112226
rect 5694 112170 5762 112226
rect 5818 112170 5886 112226
rect 5942 112170 6038 112226
rect 5418 112102 6038 112170
rect 5418 112046 5514 112102
rect 5570 112046 5638 112102
rect 5694 112046 5762 112102
rect 5818 112046 5886 112102
rect 5942 112046 6038 112102
rect 5418 111978 6038 112046
rect 5418 111922 5514 111978
rect 5570 111922 5638 111978
rect 5694 111922 5762 111978
rect 5818 111922 5886 111978
rect 5942 111922 6038 111978
rect -956 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 -336 94350
rect -956 94226 -336 94294
rect -956 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 -336 94226
rect -956 94102 -336 94170
rect -956 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 -336 94102
rect -956 93978 -336 94046
rect -956 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 -336 93978
rect -956 76350 -336 93922
rect 5418 94350 6038 111922
rect 12448 112350 12768 112384
rect 12448 112294 12518 112350
rect 12574 112294 12642 112350
rect 12698 112294 12768 112350
rect 12448 112226 12768 112294
rect 12448 112170 12518 112226
rect 12574 112170 12642 112226
rect 12698 112170 12768 112226
rect 12448 112102 12768 112170
rect 12448 112046 12518 112102
rect 12574 112046 12642 112102
rect 12698 112046 12768 112102
rect 12448 111978 12768 112046
rect 12448 111922 12518 111978
rect 12574 111922 12642 111978
rect 12698 111922 12768 111978
rect 12448 111888 12768 111922
rect 43168 112350 43488 112384
rect 43168 112294 43238 112350
rect 43294 112294 43362 112350
rect 43418 112294 43488 112350
rect 43168 112226 43488 112294
rect 43168 112170 43238 112226
rect 43294 112170 43362 112226
rect 43418 112170 43488 112226
rect 43168 112102 43488 112170
rect 43168 112046 43238 112102
rect 43294 112046 43362 112102
rect 43418 112046 43488 112102
rect 43168 111978 43488 112046
rect 43168 111922 43238 111978
rect 43294 111922 43362 111978
rect 43418 111922 43488 111978
rect 43168 111888 43488 111922
rect 73888 112350 74208 112384
rect 73888 112294 73958 112350
rect 74014 112294 74082 112350
rect 74138 112294 74208 112350
rect 73888 112226 74208 112294
rect 73888 112170 73958 112226
rect 74014 112170 74082 112226
rect 74138 112170 74208 112226
rect 73888 112102 74208 112170
rect 73888 112046 73958 112102
rect 74014 112046 74082 112102
rect 74138 112046 74208 112102
rect 73888 111978 74208 112046
rect 73888 111922 73958 111978
rect 74014 111922 74082 111978
rect 74138 111922 74208 111978
rect 73888 111888 74208 111922
rect 104608 112350 104928 112384
rect 104608 112294 104678 112350
rect 104734 112294 104802 112350
rect 104858 112294 104928 112350
rect 104608 112226 104928 112294
rect 104608 112170 104678 112226
rect 104734 112170 104802 112226
rect 104858 112170 104928 112226
rect 104608 112102 104928 112170
rect 104608 112046 104678 112102
rect 104734 112046 104802 112102
rect 104858 112046 104928 112102
rect 104608 111978 104928 112046
rect 104608 111922 104678 111978
rect 104734 111922 104802 111978
rect 104858 111922 104928 111978
rect 104608 111888 104928 111922
rect 135328 112350 135648 112384
rect 135328 112294 135398 112350
rect 135454 112294 135522 112350
rect 135578 112294 135648 112350
rect 135328 112226 135648 112294
rect 135328 112170 135398 112226
rect 135454 112170 135522 112226
rect 135578 112170 135648 112226
rect 135328 112102 135648 112170
rect 135328 112046 135398 112102
rect 135454 112046 135522 112102
rect 135578 112046 135648 112102
rect 135328 111978 135648 112046
rect 135328 111922 135398 111978
rect 135454 111922 135522 111978
rect 135578 111922 135648 111978
rect 135328 111888 135648 111922
rect 166048 112350 166368 112384
rect 166048 112294 166118 112350
rect 166174 112294 166242 112350
rect 166298 112294 166368 112350
rect 166048 112226 166368 112294
rect 166048 112170 166118 112226
rect 166174 112170 166242 112226
rect 166298 112170 166368 112226
rect 166048 112102 166368 112170
rect 166048 112046 166118 112102
rect 166174 112046 166242 112102
rect 166298 112046 166368 112102
rect 166048 111978 166368 112046
rect 166048 111922 166118 111978
rect 166174 111922 166242 111978
rect 166298 111922 166368 111978
rect 166048 111888 166368 111922
rect 196768 112350 197088 112384
rect 196768 112294 196838 112350
rect 196894 112294 196962 112350
rect 197018 112294 197088 112350
rect 196768 112226 197088 112294
rect 196768 112170 196838 112226
rect 196894 112170 196962 112226
rect 197018 112170 197088 112226
rect 196768 112102 197088 112170
rect 196768 112046 196838 112102
rect 196894 112046 196962 112102
rect 197018 112046 197088 112102
rect 196768 111978 197088 112046
rect 196768 111922 196838 111978
rect 196894 111922 196962 111978
rect 197018 111922 197088 111978
rect 196768 111888 197088 111922
rect 227488 112350 227808 112384
rect 227488 112294 227558 112350
rect 227614 112294 227682 112350
rect 227738 112294 227808 112350
rect 227488 112226 227808 112294
rect 227488 112170 227558 112226
rect 227614 112170 227682 112226
rect 227738 112170 227808 112226
rect 227488 112102 227808 112170
rect 227488 112046 227558 112102
rect 227614 112046 227682 112102
rect 227738 112046 227808 112102
rect 227488 111978 227808 112046
rect 227488 111922 227558 111978
rect 227614 111922 227682 111978
rect 227738 111922 227808 111978
rect 227488 111888 227808 111922
rect 258208 112350 258528 112384
rect 258208 112294 258278 112350
rect 258334 112294 258402 112350
rect 258458 112294 258528 112350
rect 258208 112226 258528 112294
rect 258208 112170 258278 112226
rect 258334 112170 258402 112226
rect 258458 112170 258528 112226
rect 258208 112102 258528 112170
rect 258208 112046 258278 112102
rect 258334 112046 258402 112102
rect 258458 112046 258528 112102
rect 258208 111978 258528 112046
rect 258208 111922 258278 111978
rect 258334 111922 258402 111978
rect 258458 111922 258528 111978
rect 258208 111888 258528 111922
rect 288928 112350 289248 112384
rect 288928 112294 288998 112350
rect 289054 112294 289122 112350
rect 289178 112294 289248 112350
rect 288928 112226 289248 112294
rect 288928 112170 288998 112226
rect 289054 112170 289122 112226
rect 289178 112170 289248 112226
rect 288928 112102 289248 112170
rect 288928 112046 288998 112102
rect 289054 112046 289122 112102
rect 289178 112046 289248 112102
rect 288928 111978 289248 112046
rect 288928 111922 288998 111978
rect 289054 111922 289122 111978
rect 289178 111922 289248 111978
rect 288928 111888 289248 111922
rect 319648 112350 319968 112384
rect 319648 112294 319718 112350
rect 319774 112294 319842 112350
rect 319898 112294 319968 112350
rect 319648 112226 319968 112294
rect 319648 112170 319718 112226
rect 319774 112170 319842 112226
rect 319898 112170 319968 112226
rect 319648 112102 319968 112170
rect 319648 112046 319718 112102
rect 319774 112046 319842 112102
rect 319898 112046 319968 112102
rect 319648 111978 319968 112046
rect 319648 111922 319718 111978
rect 319774 111922 319842 111978
rect 319898 111922 319968 111978
rect 319648 111888 319968 111922
rect 350368 112350 350688 112384
rect 350368 112294 350438 112350
rect 350494 112294 350562 112350
rect 350618 112294 350688 112350
rect 350368 112226 350688 112294
rect 350368 112170 350438 112226
rect 350494 112170 350562 112226
rect 350618 112170 350688 112226
rect 350368 112102 350688 112170
rect 350368 112046 350438 112102
rect 350494 112046 350562 112102
rect 350618 112046 350688 112102
rect 350368 111978 350688 112046
rect 350368 111922 350438 111978
rect 350494 111922 350562 111978
rect 350618 111922 350688 111978
rect 350368 111888 350688 111922
rect 381088 112350 381408 112384
rect 381088 112294 381158 112350
rect 381214 112294 381282 112350
rect 381338 112294 381408 112350
rect 381088 112226 381408 112294
rect 381088 112170 381158 112226
rect 381214 112170 381282 112226
rect 381338 112170 381408 112226
rect 381088 112102 381408 112170
rect 381088 112046 381158 112102
rect 381214 112046 381282 112102
rect 381338 112046 381408 112102
rect 381088 111978 381408 112046
rect 381088 111922 381158 111978
rect 381214 111922 381282 111978
rect 381338 111922 381408 111978
rect 381088 111888 381408 111922
rect 411808 112350 412128 112384
rect 411808 112294 411878 112350
rect 411934 112294 412002 112350
rect 412058 112294 412128 112350
rect 411808 112226 412128 112294
rect 411808 112170 411878 112226
rect 411934 112170 412002 112226
rect 412058 112170 412128 112226
rect 411808 112102 412128 112170
rect 411808 112046 411878 112102
rect 411934 112046 412002 112102
rect 412058 112046 412128 112102
rect 411808 111978 412128 112046
rect 411808 111922 411878 111978
rect 411934 111922 412002 111978
rect 412058 111922 412128 111978
rect 411808 111888 412128 111922
rect 442528 112350 442848 112384
rect 442528 112294 442598 112350
rect 442654 112294 442722 112350
rect 442778 112294 442848 112350
rect 442528 112226 442848 112294
rect 442528 112170 442598 112226
rect 442654 112170 442722 112226
rect 442778 112170 442848 112226
rect 442528 112102 442848 112170
rect 442528 112046 442598 112102
rect 442654 112046 442722 112102
rect 442778 112046 442848 112102
rect 442528 111978 442848 112046
rect 442528 111922 442598 111978
rect 442654 111922 442722 111978
rect 442778 111922 442848 111978
rect 442528 111888 442848 111922
rect 473248 112350 473568 112384
rect 473248 112294 473318 112350
rect 473374 112294 473442 112350
rect 473498 112294 473568 112350
rect 473248 112226 473568 112294
rect 473248 112170 473318 112226
rect 473374 112170 473442 112226
rect 473498 112170 473568 112226
rect 473248 112102 473568 112170
rect 473248 112046 473318 112102
rect 473374 112046 473442 112102
rect 473498 112046 473568 112102
rect 473248 111978 473568 112046
rect 473248 111922 473318 111978
rect 473374 111922 473442 111978
rect 473498 111922 473568 111978
rect 473248 111888 473568 111922
rect 503968 112350 504288 112384
rect 503968 112294 504038 112350
rect 504094 112294 504162 112350
rect 504218 112294 504288 112350
rect 503968 112226 504288 112294
rect 503968 112170 504038 112226
rect 504094 112170 504162 112226
rect 504218 112170 504288 112226
rect 503968 112102 504288 112170
rect 503968 112046 504038 112102
rect 504094 112046 504162 112102
rect 504218 112046 504288 112102
rect 503968 111978 504288 112046
rect 503968 111922 504038 111978
rect 504094 111922 504162 111978
rect 504218 111922 504288 111978
rect 503968 111888 504288 111922
rect 534688 112350 535008 112384
rect 534688 112294 534758 112350
rect 534814 112294 534882 112350
rect 534938 112294 535008 112350
rect 534688 112226 535008 112294
rect 534688 112170 534758 112226
rect 534814 112170 534882 112226
rect 534938 112170 535008 112226
rect 534688 112102 535008 112170
rect 534688 112046 534758 112102
rect 534814 112046 534882 112102
rect 534938 112046 535008 112102
rect 534688 111978 535008 112046
rect 534688 111922 534758 111978
rect 534814 111922 534882 111978
rect 534938 111922 535008 111978
rect 534688 111888 535008 111922
rect 565408 112350 565728 112384
rect 565408 112294 565478 112350
rect 565534 112294 565602 112350
rect 565658 112294 565728 112350
rect 565408 112226 565728 112294
rect 565408 112170 565478 112226
rect 565534 112170 565602 112226
rect 565658 112170 565728 112226
rect 565408 112102 565728 112170
rect 565408 112046 565478 112102
rect 565534 112046 565602 112102
rect 565658 112046 565728 112102
rect 565408 111978 565728 112046
rect 565408 111922 565478 111978
rect 565534 111922 565602 111978
rect 565658 111922 565728 111978
rect 565408 111888 565728 111922
rect 589098 112350 589718 129922
rect 590492 139300 590548 139310
rect 590492 124740 590548 139244
rect 592818 136350 593438 153922
rect 592818 136294 592914 136350
rect 592970 136294 593038 136350
rect 593094 136294 593162 136350
rect 593218 136294 593286 136350
rect 593342 136294 593438 136350
rect 592818 136226 593438 136294
rect 592818 136170 592914 136226
rect 592970 136170 593038 136226
rect 593094 136170 593162 136226
rect 593218 136170 593286 136226
rect 593342 136170 593438 136226
rect 592818 136102 593438 136170
rect 592818 136046 592914 136102
rect 592970 136046 593038 136102
rect 593094 136046 593162 136102
rect 593218 136046 593286 136102
rect 593342 136046 593438 136102
rect 592818 135978 593438 136046
rect 592818 135922 592914 135978
rect 592970 135922 593038 135978
rect 593094 135922 593162 135978
rect 593218 135922 593286 135978
rect 593342 135922 593438 135978
rect 590492 124674 590548 124684
rect 590604 126084 590660 126094
rect 590604 113988 590660 126028
rect 590604 113922 590660 113932
rect 592818 118350 593438 135922
rect 592818 118294 592914 118350
rect 592970 118294 593038 118350
rect 593094 118294 593162 118350
rect 593218 118294 593286 118350
rect 593342 118294 593438 118350
rect 592818 118226 593438 118294
rect 592818 118170 592914 118226
rect 592970 118170 593038 118226
rect 593094 118170 593162 118226
rect 593218 118170 593286 118226
rect 593342 118170 593438 118226
rect 592818 118102 593438 118170
rect 592818 118046 592914 118102
rect 592970 118046 593038 118102
rect 593094 118046 593162 118102
rect 593218 118046 593286 118102
rect 593342 118046 593438 118102
rect 592818 117978 593438 118046
rect 592818 117922 592914 117978
rect 592970 117922 593038 117978
rect 593094 117922 593162 117978
rect 593218 117922 593286 117978
rect 593342 117922 593438 117978
rect 589098 112294 589194 112350
rect 589250 112294 589318 112350
rect 589374 112294 589442 112350
rect 589498 112294 589566 112350
rect 589622 112294 589718 112350
rect 589098 112226 589718 112294
rect 589098 112170 589194 112226
rect 589250 112170 589318 112226
rect 589374 112170 589442 112226
rect 589498 112170 589566 112226
rect 589622 112170 589718 112226
rect 589098 112102 589718 112170
rect 589098 112046 589194 112102
rect 589250 112046 589318 112102
rect 589374 112046 589442 112102
rect 589498 112046 589566 112102
rect 589622 112046 589718 112102
rect 589098 111978 589718 112046
rect 589098 111922 589194 111978
rect 589250 111922 589318 111978
rect 589374 111922 589442 111978
rect 589498 111922 589566 111978
rect 589622 111922 589718 111978
rect 5418 94294 5514 94350
rect 5570 94294 5638 94350
rect 5694 94294 5762 94350
rect 5818 94294 5886 94350
rect 5942 94294 6038 94350
rect 5418 94226 6038 94294
rect 5418 94170 5514 94226
rect 5570 94170 5638 94226
rect 5694 94170 5762 94226
rect 5818 94170 5886 94226
rect 5942 94170 6038 94226
rect 5418 94102 6038 94170
rect 5418 94046 5514 94102
rect 5570 94046 5638 94102
rect 5694 94046 5762 94102
rect 5818 94046 5886 94102
rect 5942 94046 6038 94102
rect 5418 93978 6038 94046
rect 5418 93922 5514 93978
rect 5570 93922 5638 93978
rect 5694 93922 5762 93978
rect 5818 93922 5886 93978
rect 5942 93922 6038 93978
rect 4172 93268 4228 93278
rect 4172 80836 4228 93212
rect 4172 80770 4228 80780
rect -956 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 -336 76350
rect -956 76226 -336 76294
rect -956 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 -336 76226
rect -956 76102 -336 76170
rect -956 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 -336 76102
rect -956 75978 -336 76046
rect -956 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 -336 75978
rect -956 58350 -336 75922
rect 4172 79156 4228 79166
rect 4172 70308 4228 79100
rect 4172 70242 4228 70252
rect 5418 76350 6038 93922
rect 6188 107380 6244 107390
rect 6188 91364 6244 107324
rect 27808 100350 28128 100384
rect 27808 100294 27878 100350
rect 27934 100294 28002 100350
rect 28058 100294 28128 100350
rect 27808 100226 28128 100294
rect 27808 100170 27878 100226
rect 27934 100170 28002 100226
rect 28058 100170 28128 100226
rect 27808 100102 28128 100170
rect 27808 100046 27878 100102
rect 27934 100046 28002 100102
rect 28058 100046 28128 100102
rect 27808 99978 28128 100046
rect 27808 99922 27878 99978
rect 27934 99922 28002 99978
rect 28058 99922 28128 99978
rect 27808 99888 28128 99922
rect 58528 100350 58848 100384
rect 58528 100294 58598 100350
rect 58654 100294 58722 100350
rect 58778 100294 58848 100350
rect 58528 100226 58848 100294
rect 58528 100170 58598 100226
rect 58654 100170 58722 100226
rect 58778 100170 58848 100226
rect 58528 100102 58848 100170
rect 58528 100046 58598 100102
rect 58654 100046 58722 100102
rect 58778 100046 58848 100102
rect 58528 99978 58848 100046
rect 58528 99922 58598 99978
rect 58654 99922 58722 99978
rect 58778 99922 58848 99978
rect 58528 99888 58848 99922
rect 89248 100350 89568 100384
rect 89248 100294 89318 100350
rect 89374 100294 89442 100350
rect 89498 100294 89568 100350
rect 89248 100226 89568 100294
rect 89248 100170 89318 100226
rect 89374 100170 89442 100226
rect 89498 100170 89568 100226
rect 89248 100102 89568 100170
rect 89248 100046 89318 100102
rect 89374 100046 89442 100102
rect 89498 100046 89568 100102
rect 89248 99978 89568 100046
rect 89248 99922 89318 99978
rect 89374 99922 89442 99978
rect 89498 99922 89568 99978
rect 89248 99888 89568 99922
rect 119968 100350 120288 100384
rect 119968 100294 120038 100350
rect 120094 100294 120162 100350
rect 120218 100294 120288 100350
rect 119968 100226 120288 100294
rect 119968 100170 120038 100226
rect 120094 100170 120162 100226
rect 120218 100170 120288 100226
rect 119968 100102 120288 100170
rect 119968 100046 120038 100102
rect 120094 100046 120162 100102
rect 120218 100046 120288 100102
rect 119968 99978 120288 100046
rect 119968 99922 120038 99978
rect 120094 99922 120162 99978
rect 120218 99922 120288 99978
rect 119968 99888 120288 99922
rect 150688 100350 151008 100384
rect 150688 100294 150758 100350
rect 150814 100294 150882 100350
rect 150938 100294 151008 100350
rect 150688 100226 151008 100294
rect 150688 100170 150758 100226
rect 150814 100170 150882 100226
rect 150938 100170 151008 100226
rect 150688 100102 151008 100170
rect 150688 100046 150758 100102
rect 150814 100046 150882 100102
rect 150938 100046 151008 100102
rect 150688 99978 151008 100046
rect 150688 99922 150758 99978
rect 150814 99922 150882 99978
rect 150938 99922 151008 99978
rect 150688 99888 151008 99922
rect 181408 100350 181728 100384
rect 181408 100294 181478 100350
rect 181534 100294 181602 100350
rect 181658 100294 181728 100350
rect 181408 100226 181728 100294
rect 181408 100170 181478 100226
rect 181534 100170 181602 100226
rect 181658 100170 181728 100226
rect 181408 100102 181728 100170
rect 181408 100046 181478 100102
rect 181534 100046 181602 100102
rect 181658 100046 181728 100102
rect 181408 99978 181728 100046
rect 181408 99922 181478 99978
rect 181534 99922 181602 99978
rect 181658 99922 181728 99978
rect 181408 99888 181728 99922
rect 212128 100350 212448 100384
rect 212128 100294 212198 100350
rect 212254 100294 212322 100350
rect 212378 100294 212448 100350
rect 212128 100226 212448 100294
rect 212128 100170 212198 100226
rect 212254 100170 212322 100226
rect 212378 100170 212448 100226
rect 212128 100102 212448 100170
rect 212128 100046 212198 100102
rect 212254 100046 212322 100102
rect 212378 100046 212448 100102
rect 212128 99978 212448 100046
rect 212128 99922 212198 99978
rect 212254 99922 212322 99978
rect 212378 99922 212448 99978
rect 212128 99888 212448 99922
rect 242848 100350 243168 100384
rect 242848 100294 242918 100350
rect 242974 100294 243042 100350
rect 243098 100294 243168 100350
rect 242848 100226 243168 100294
rect 242848 100170 242918 100226
rect 242974 100170 243042 100226
rect 243098 100170 243168 100226
rect 242848 100102 243168 100170
rect 242848 100046 242918 100102
rect 242974 100046 243042 100102
rect 243098 100046 243168 100102
rect 242848 99978 243168 100046
rect 242848 99922 242918 99978
rect 242974 99922 243042 99978
rect 243098 99922 243168 99978
rect 242848 99888 243168 99922
rect 273568 100350 273888 100384
rect 273568 100294 273638 100350
rect 273694 100294 273762 100350
rect 273818 100294 273888 100350
rect 273568 100226 273888 100294
rect 273568 100170 273638 100226
rect 273694 100170 273762 100226
rect 273818 100170 273888 100226
rect 273568 100102 273888 100170
rect 273568 100046 273638 100102
rect 273694 100046 273762 100102
rect 273818 100046 273888 100102
rect 273568 99978 273888 100046
rect 273568 99922 273638 99978
rect 273694 99922 273762 99978
rect 273818 99922 273888 99978
rect 273568 99888 273888 99922
rect 304288 100350 304608 100384
rect 304288 100294 304358 100350
rect 304414 100294 304482 100350
rect 304538 100294 304608 100350
rect 304288 100226 304608 100294
rect 304288 100170 304358 100226
rect 304414 100170 304482 100226
rect 304538 100170 304608 100226
rect 304288 100102 304608 100170
rect 304288 100046 304358 100102
rect 304414 100046 304482 100102
rect 304538 100046 304608 100102
rect 304288 99978 304608 100046
rect 304288 99922 304358 99978
rect 304414 99922 304482 99978
rect 304538 99922 304608 99978
rect 304288 99888 304608 99922
rect 335008 100350 335328 100384
rect 335008 100294 335078 100350
rect 335134 100294 335202 100350
rect 335258 100294 335328 100350
rect 335008 100226 335328 100294
rect 335008 100170 335078 100226
rect 335134 100170 335202 100226
rect 335258 100170 335328 100226
rect 335008 100102 335328 100170
rect 335008 100046 335078 100102
rect 335134 100046 335202 100102
rect 335258 100046 335328 100102
rect 335008 99978 335328 100046
rect 335008 99922 335078 99978
rect 335134 99922 335202 99978
rect 335258 99922 335328 99978
rect 335008 99888 335328 99922
rect 365728 100350 366048 100384
rect 365728 100294 365798 100350
rect 365854 100294 365922 100350
rect 365978 100294 366048 100350
rect 365728 100226 366048 100294
rect 365728 100170 365798 100226
rect 365854 100170 365922 100226
rect 365978 100170 366048 100226
rect 365728 100102 366048 100170
rect 365728 100046 365798 100102
rect 365854 100046 365922 100102
rect 365978 100046 366048 100102
rect 365728 99978 366048 100046
rect 365728 99922 365798 99978
rect 365854 99922 365922 99978
rect 365978 99922 366048 99978
rect 365728 99888 366048 99922
rect 396448 100350 396768 100384
rect 396448 100294 396518 100350
rect 396574 100294 396642 100350
rect 396698 100294 396768 100350
rect 396448 100226 396768 100294
rect 396448 100170 396518 100226
rect 396574 100170 396642 100226
rect 396698 100170 396768 100226
rect 396448 100102 396768 100170
rect 396448 100046 396518 100102
rect 396574 100046 396642 100102
rect 396698 100046 396768 100102
rect 396448 99978 396768 100046
rect 396448 99922 396518 99978
rect 396574 99922 396642 99978
rect 396698 99922 396768 99978
rect 396448 99888 396768 99922
rect 427168 100350 427488 100384
rect 427168 100294 427238 100350
rect 427294 100294 427362 100350
rect 427418 100294 427488 100350
rect 427168 100226 427488 100294
rect 427168 100170 427238 100226
rect 427294 100170 427362 100226
rect 427418 100170 427488 100226
rect 427168 100102 427488 100170
rect 427168 100046 427238 100102
rect 427294 100046 427362 100102
rect 427418 100046 427488 100102
rect 427168 99978 427488 100046
rect 427168 99922 427238 99978
rect 427294 99922 427362 99978
rect 427418 99922 427488 99978
rect 427168 99888 427488 99922
rect 457888 100350 458208 100384
rect 457888 100294 457958 100350
rect 458014 100294 458082 100350
rect 458138 100294 458208 100350
rect 457888 100226 458208 100294
rect 457888 100170 457958 100226
rect 458014 100170 458082 100226
rect 458138 100170 458208 100226
rect 457888 100102 458208 100170
rect 457888 100046 457958 100102
rect 458014 100046 458082 100102
rect 458138 100046 458208 100102
rect 457888 99978 458208 100046
rect 457888 99922 457958 99978
rect 458014 99922 458082 99978
rect 458138 99922 458208 99978
rect 457888 99888 458208 99922
rect 488608 100350 488928 100384
rect 488608 100294 488678 100350
rect 488734 100294 488802 100350
rect 488858 100294 488928 100350
rect 488608 100226 488928 100294
rect 488608 100170 488678 100226
rect 488734 100170 488802 100226
rect 488858 100170 488928 100226
rect 488608 100102 488928 100170
rect 488608 100046 488678 100102
rect 488734 100046 488802 100102
rect 488858 100046 488928 100102
rect 488608 99978 488928 100046
rect 488608 99922 488678 99978
rect 488734 99922 488802 99978
rect 488858 99922 488928 99978
rect 488608 99888 488928 99922
rect 519328 100350 519648 100384
rect 519328 100294 519398 100350
rect 519454 100294 519522 100350
rect 519578 100294 519648 100350
rect 519328 100226 519648 100294
rect 519328 100170 519398 100226
rect 519454 100170 519522 100226
rect 519578 100170 519648 100226
rect 519328 100102 519648 100170
rect 519328 100046 519398 100102
rect 519454 100046 519522 100102
rect 519578 100046 519648 100102
rect 519328 99978 519648 100046
rect 519328 99922 519398 99978
rect 519454 99922 519522 99978
rect 519578 99922 519648 99978
rect 519328 99888 519648 99922
rect 550048 100350 550368 100384
rect 550048 100294 550118 100350
rect 550174 100294 550242 100350
rect 550298 100294 550368 100350
rect 550048 100226 550368 100294
rect 550048 100170 550118 100226
rect 550174 100170 550242 100226
rect 550298 100170 550368 100226
rect 550048 100102 550368 100170
rect 550048 100046 550118 100102
rect 550174 100046 550242 100102
rect 550298 100046 550368 100102
rect 550048 99978 550368 100046
rect 550048 99922 550118 99978
rect 550174 99922 550242 99978
rect 550298 99922 550368 99978
rect 550048 99888 550368 99922
rect 587132 99652 587188 99662
rect 12448 94350 12768 94384
rect 12448 94294 12518 94350
rect 12574 94294 12642 94350
rect 12698 94294 12768 94350
rect 12448 94226 12768 94294
rect 12448 94170 12518 94226
rect 12574 94170 12642 94226
rect 12698 94170 12768 94226
rect 12448 94102 12768 94170
rect 12448 94046 12518 94102
rect 12574 94046 12642 94102
rect 12698 94046 12768 94102
rect 12448 93978 12768 94046
rect 12448 93922 12518 93978
rect 12574 93922 12642 93978
rect 12698 93922 12768 93978
rect 12448 93888 12768 93922
rect 43168 94350 43488 94384
rect 43168 94294 43238 94350
rect 43294 94294 43362 94350
rect 43418 94294 43488 94350
rect 43168 94226 43488 94294
rect 43168 94170 43238 94226
rect 43294 94170 43362 94226
rect 43418 94170 43488 94226
rect 43168 94102 43488 94170
rect 43168 94046 43238 94102
rect 43294 94046 43362 94102
rect 43418 94046 43488 94102
rect 43168 93978 43488 94046
rect 43168 93922 43238 93978
rect 43294 93922 43362 93978
rect 43418 93922 43488 93978
rect 43168 93888 43488 93922
rect 73888 94350 74208 94384
rect 73888 94294 73958 94350
rect 74014 94294 74082 94350
rect 74138 94294 74208 94350
rect 73888 94226 74208 94294
rect 73888 94170 73958 94226
rect 74014 94170 74082 94226
rect 74138 94170 74208 94226
rect 73888 94102 74208 94170
rect 73888 94046 73958 94102
rect 74014 94046 74082 94102
rect 74138 94046 74208 94102
rect 73888 93978 74208 94046
rect 73888 93922 73958 93978
rect 74014 93922 74082 93978
rect 74138 93922 74208 93978
rect 73888 93888 74208 93922
rect 104608 94350 104928 94384
rect 104608 94294 104678 94350
rect 104734 94294 104802 94350
rect 104858 94294 104928 94350
rect 104608 94226 104928 94294
rect 104608 94170 104678 94226
rect 104734 94170 104802 94226
rect 104858 94170 104928 94226
rect 104608 94102 104928 94170
rect 104608 94046 104678 94102
rect 104734 94046 104802 94102
rect 104858 94046 104928 94102
rect 104608 93978 104928 94046
rect 104608 93922 104678 93978
rect 104734 93922 104802 93978
rect 104858 93922 104928 93978
rect 104608 93888 104928 93922
rect 135328 94350 135648 94384
rect 135328 94294 135398 94350
rect 135454 94294 135522 94350
rect 135578 94294 135648 94350
rect 135328 94226 135648 94294
rect 135328 94170 135398 94226
rect 135454 94170 135522 94226
rect 135578 94170 135648 94226
rect 135328 94102 135648 94170
rect 135328 94046 135398 94102
rect 135454 94046 135522 94102
rect 135578 94046 135648 94102
rect 135328 93978 135648 94046
rect 135328 93922 135398 93978
rect 135454 93922 135522 93978
rect 135578 93922 135648 93978
rect 135328 93888 135648 93922
rect 166048 94350 166368 94384
rect 166048 94294 166118 94350
rect 166174 94294 166242 94350
rect 166298 94294 166368 94350
rect 166048 94226 166368 94294
rect 166048 94170 166118 94226
rect 166174 94170 166242 94226
rect 166298 94170 166368 94226
rect 166048 94102 166368 94170
rect 166048 94046 166118 94102
rect 166174 94046 166242 94102
rect 166298 94046 166368 94102
rect 166048 93978 166368 94046
rect 166048 93922 166118 93978
rect 166174 93922 166242 93978
rect 166298 93922 166368 93978
rect 166048 93888 166368 93922
rect 196768 94350 197088 94384
rect 196768 94294 196838 94350
rect 196894 94294 196962 94350
rect 197018 94294 197088 94350
rect 196768 94226 197088 94294
rect 196768 94170 196838 94226
rect 196894 94170 196962 94226
rect 197018 94170 197088 94226
rect 196768 94102 197088 94170
rect 196768 94046 196838 94102
rect 196894 94046 196962 94102
rect 197018 94046 197088 94102
rect 196768 93978 197088 94046
rect 196768 93922 196838 93978
rect 196894 93922 196962 93978
rect 197018 93922 197088 93978
rect 196768 93888 197088 93922
rect 227488 94350 227808 94384
rect 227488 94294 227558 94350
rect 227614 94294 227682 94350
rect 227738 94294 227808 94350
rect 227488 94226 227808 94294
rect 227488 94170 227558 94226
rect 227614 94170 227682 94226
rect 227738 94170 227808 94226
rect 227488 94102 227808 94170
rect 227488 94046 227558 94102
rect 227614 94046 227682 94102
rect 227738 94046 227808 94102
rect 227488 93978 227808 94046
rect 227488 93922 227558 93978
rect 227614 93922 227682 93978
rect 227738 93922 227808 93978
rect 227488 93888 227808 93922
rect 258208 94350 258528 94384
rect 258208 94294 258278 94350
rect 258334 94294 258402 94350
rect 258458 94294 258528 94350
rect 258208 94226 258528 94294
rect 258208 94170 258278 94226
rect 258334 94170 258402 94226
rect 258458 94170 258528 94226
rect 258208 94102 258528 94170
rect 258208 94046 258278 94102
rect 258334 94046 258402 94102
rect 258458 94046 258528 94102
rect 258208 93978 258528 94046
rect 258208 93922 258278 93978
rect 258334 93922 258402 93978
rect 258458 93922 258528 93978
rect 258208 93888 258528 93922
rect 288928 94350 289248 94384
rect 288928 94294 288998 94350
rect 289054 94294 289122 94350
rect 289178 94294 289248 94350
rect 288928 94226 289248 94294
rect 288928 94170 288998 94226
rect 289054 94170 289122 94226
rect 289178 94170 289248 94226
rect 288928 94102 289248 94170
rect 288928 94046 288998 94102
rect 289054 94046 289122 94102
rect 289178 94046 289248 94102
rect 288928 93978 289248 94046
rect 288928 93922 288998 93978
rect 289054 93922 289122 93978
rect 289178 93922 289248 93978
rect 288928 93888 289248 93922
rect 319648 94350 319968 94384
rect 319648 94294 319718 94350
rect 319774 94294 319842 94350
rect 319898 94294 319968 94350
rect 319648 94226 319968 94294
rect 319648 94170 319718 94226
rect 319774 94170 319842 94226
rect 319898 94170 319968 94226
rect 319648 94102 319968 94170
rect 319648 94046 319718 94102
rect 319774 94046 319842 94102
rect 319898 94046 319968 94102
rect 319648 93978 319968 94046
rect 319648 93922 319718 93978
rect 319774 93922 319842 93978
rect 319898 93922 319968 93978
rect 319648 93888 319968 93922
rect 350368 94350 350688 94384
rect 350368 94294 350438 94350
rect 350494 94294 350562 94350
rect 350618 94294 350688 94350
rect 350368 94226 350688 94294
rect 350368 94170 350438 94226
rect 350494 94170 350562 94226
rect 350618 94170 350688 94226
rect 350368 94102 350688 94170
rect 350368 94046 350438 94102
rect 350494 94046 350562 94102
rect 350618 94046 350688 94102
rect 350368 93978 350688 94046
rect 350368 93922 350438 93978
rect 350494 93922 350562 93978
rect 350618 93922 350688 93978
rect 350368 93888 350688 93922
rect 381088 94350 381408 94384
rect 381088 94294 381158 94350
rect 381214 94294 381282 94350
rect 381338 94294 381408 94350
rect 381088 94226 381408 94294
rect 381088 94170 381158 94226
rect 381214 94170 381282 94226
rect 381338 94170 381408 94226
rect 381088 94102 381408 94170
rect 381088 94046 381158 94102
rect 381214 94046 381282 94102
rect 381338 94046 381408 94102
rect 381088 93978 381408 94046
rect 381088 93922 381158 93978
rect 381214 93922 381282 93978
rect 381338 93922 381408 93978
rect 381088 93888 381408 93922
rect 411808 94350 412128 94384
rect 411808 94294 411878 94350
rect 411934 94294 412002 94350
rect 412058 94294 412128 94350
rect 411808 94226 412128 94294
rect 411808 94170 411878 94226
rect 411934 94170 412002 94226
rect 412058 94170 412128 94226
rect 411808 94102 412128 94170
rect 411808 94046 411878 94102
rect 411934 94046 412002 94102
rect 412058 94046 412128 94102
rect 411808 93978 412128 94046
rect 411808 93922 411878 93978
rect 411934 93922 412002 93978
rect 412058 93922 412128 93978
rect 411808 93888 412128 93922
rect 442528 94350 442848 94384
rect 442528 94294 442598 94350
rect 442654 94294 442722 94350
rect 442778 94294 442848 94350
rect 442528 94226 442848 94294
rect 442528 94170 442598 94226
rect 442654 94170 442722 94226
rect 442778 94170 442848 94226
rect 442528 94102 442848 94170
rect 442528 94046 442598 94102
rect 442654 94046 442722 94102
rect 442778 94046 442848 94102
rect 442528 93978 442848 94046
rect 442528 93922 442598 93978
rect 442654 93922 442722 93978
rect 442778 93922 442848 93978
rect 442528 93888 442848 93922
rect 473248 94350 473568 94384
rect 473248 94294 473318 94350
rect 473374 94294 473442 94350
rect 473498 94294 473568 94350
rect 473248 94226 473568 94294
rect 473248 94170 473318 94226
rect 473374 94170 473442 94226
rect 473498 94170 473568 94226
rect 473248 94102 473568 94170
rect 473248 94046 473318 94102
rect 473374 94046 473442 94102
rect 473498 94046 473568 94102
rect 473248 93978 473568 94046
rect 473248 93922 473318 93978
rect 473374 93922 473442 93978
rect 473498 93922 473568 93978
rect 473248 93888 473568 93922
rect 503968 94350 504288 94384
rect 503968 94294 504038 94350
rect 504094 94294 504162 94350
rect 504218 94294 504288 94350
rect 503968 94226 504288 94294
rect 503968 94170 504038 94226
rect 504094 94170 504162 94226
rect 504218 94170 504288 94226
rect 503968 94102 504288 94170
rect 503968 94046 504038 94102
rect 504094 94046 504162 94102
rect 504218 94046 504288 94102
rect 503968 93978 504288 94046
rect 503968 93922 504038 93978
rect 504094 93922 504162 93978
rect 504218 93922 504288 93978
rect 503968 93888 504288 93922
rect 534688 94350 535008 94384
rect 534688 94294 534758 94350
rect 534814 94294 534882 94350
rect 534938 94294 535008 94350
rect 534688 94226 535008 94294
rect 534688 94170 534758 94226
rect 534814 94170 534882 94226
rect 534938 94170 535008 94226
rect 534688 94102 535008 94170
rect 534688 94046 534758 94102
rect 534814 94046 534882 94102
rect 534938 94046 535008 94102
rect 534688 93978 535008 94046
rect 534688 93922 534758 93978
rect 534814 93922 534882 93978
rect 534938 93922 535008 93978
rect 534688 93888 535008 93922
rect 565408 94350 565728 94384
rect 565408 94294 565478 94350
rect 565534 94294 565602 94350
rect 565658 94294 565728 94350
rect 565408 94226 565728 94294
rect 565408 94170 565478 94226
rect 565534 94170 565602 94226
rect 565658 94170 565728 94226
rect 565408 94102 565728 94170
rect 565408 94046 565478 94102
rect 565534 94046 565602 94102
rect 565658 94046 565728 94102
rect 565408 93978 565728 94046
rect 565408 93922 565478 93978
rect 565534 93922 565602 93978
rect 565658 93922 565728 93978
rect 565408 93888 565728 93922
rect 587132 92484 587188 99596
rect 587132 92418 587188 92428
rect 589098 94350 589718 111922
rect 590828 112868 590884 112878
rect 590828 103236 590884 112812
rect 590828 103170 590884 103180
rect 589098 94294 589194 94350
rect 589250 94294 589318 94350
rect 589374 94294 589442 94350
rect 589498 94294 589566 94350
rect 589622 94294 589718 94350
rect 589098 94226 589718 94294
rect 589098 94170 589194 94226
rect 589250 94170 589318 94226
rect 589374 94170 589442 94226
rect 589498 94170 589566 94226
rect 589622 94170 589718 94226
rect 589098 94102 589718 94170
rect 589098 94046 589194 94102
rect 589250 94046 589318 94102
rect 589374 94046 589442 94102
rect 589498 94046 589566 94102
rect 589622 94046 589718 94102
rect 589098 93978 589718 94046
rect 589098 93922 589194 93978
rect 589250 93922 589318 93978
rect 589374 93922 589442 93978
rect 589498 93922 589566 93978
rect 589622 93922 589718 93978
rect 6188 91298 6244 91308
rect 27808 82350 28128 82384
rect 27808 82294 27878 82350
rect 27934 82294 28002 82350
rect 28058 82294 28128 82350
rect 27808 82226 28128 82294
rect 27808 82170 27878 82226
rect 27934 82170 28002 82226
rect 28058 82170 28128 82226
rect 27808 82102 28128 82170
rect 27808 82046 27878 82102
rect 27934 82046 28002 82102
rect 28058 82046 28128 82102
rect 27808 81978 28128 82046
rect 27808 81922 27878 81978
rect 27934 81922 28002 81978
rect 28058 81922 28128 81978
rect 27808 81888 28128 81922
rect 58528 82350 58848 82384
rect 58528 82294 58598 82350
rect 58654 82294 58722 82350
rect 58778 82294 58848 82350
rect 58528 82226 58848 82294
rect 58528 82170 58598 82226
rect 58654 82170 58722 82226
rect 58778 82170 58848 82226
rect 58528 82102 58848 82170
rect 58528 82046 58598 82102
rect 58654 82046 58722 82102
rect 58778 82046 58848 82102
rect 58528 81978 58848 82046
rect 58528 81922 58598 81978
rect 58654 81922 58722 81978
rect 58778 81922 58848 81978
rect 58528 81888 58848 81922
rect 89248 82350 89568 82384
rect 89248 82294 89318 82350
rect 89374 82294 89442 82350
rect 89498 82294 89568 82350
rect 89248 82226 89568 82294
rect 89248 82170 89318 82226
rect 89374 82170 89442 82226
rect 89498 82170 89568 82226
rect 89248 82102 89568 82170
rect 89248 82046 89318 82102
rect 89374 82046 89442 82102
rect 89498 82046 89568 82102
rect 89248 81978 89568 82046
rect 89248 81922 89318 81978
rect 89374 81922 89442 81978
rect 89498 81922 89568 81978
rect 89248 81888 89568 81922
rect 119968 82350 120288 82384
rect 119968 82294 120038 82350
rect 120094 82294 120162 82350
rect 120218 82294 120288 82350
rect 119968 82226 120288 82294
rect 119968 82170 120038 82226
rect 120094 82170 120162 82226
rect 120218 82170 120288 82226
rect 119968 82102 120288 82170
rect 119968 82046 120038 82102
rect 120094 82046 120162 82102
rect 120218 82046 120288 82102
rect 119968 81978 120288 82046
rect 119968 81922 120038 81978
rect 120094 81922 120162 81978
rect 120218 81922 120288 81978
rect 119968 81888 120288 81922
rect 150688 82350 151008 82384
rect 150688 82294 150758 82350
rect 150814 82294 150882 82350
rect 150938 82294 151008 82350
rect 150688 82226 151008 82294
rect 150688 82170 150758 82226
rect 150814 82170 150882 82226
rect 150938 82170 151008 82226
rect 150688 82102 151008 82170
rect 150688 82046 150758 82102
rect 150814 82046 150882 82102
rect 150938 82046 151008 82102
rect 150688 81978 151008 82046
rect 150688 81922 150758 81978
rect 150814 81922 150882 81978
rect 150938 81922 151008 81978
rect 150688 81888 151008 81922
rect 181408 82350 181728 82384
rect 181408 82294 181478 82350
rect 181534 82294 181602 82350
rect 181658 82294 181728 82350
rect 181408 82226 181728 82294
rect 181408 82170 181478 82226
rect 181534 82170 181602 82226
rect 181658 82170 181728 82226
rect 181408 82102 181728 82170
rect 181408 82046 181478 82102
rect 181534 82046 181602 82102
rect 181658 82046 181728 82102
rect 181408 81978 181728 82046
rect 181408 81922 181478 81978
rect 181534 81922 181602 81978
rect 181658 81922 181728 81978
rect 181408 81888 181728 81922
rect 212128 82350 212448 82384
rect 212128 82294 212198 82350
rect 212254 82294 212322 82350
rect 212378 82294 212448 82350
rect 212128 82226 212448 82294
rect 212128 82170 212198 82226
rect 212254 82170 212322 82226
rect 212378 82170 212448 82226
rect 212128 82102 212448 82170
rect 212128 82046 212198 82102
rect 212254 82046 212322 82102
rect 212378 82046 212448 82102
rect 212128 81978 212448 82046
rect 212128 81922 212198 81978
rect 212254 81922 212322 81978
rect 212378 81922 212448 81978
rect 212128 81888 212448 81922
rect 242848 82350 243168 82384
rect 242848 82294 242918 82350
rect 242974 82294 243042 82350
rect 243098 82294 243168 82350
rect 242848 82226 243168 82294
rect 242848 82170 242918 82226
rect 242974 82170 243042 82226
rect 243098 82170 243168 82226
rect 242848 82102 243168 82170
rect 242848 82046 242918 82102
rect 242974 82046 243042 82102
rect 243098 82046 243168 82102
rect 242848 81978 243168 82046
rect 242848 81922 242918 81978
rect 242974 81922 243042 81978
rect 243098 81922 243168 81978
rect 242848 81888 243168 81922
rect 273568 82350 273888 82384
rect 273568 82294 273638 82350
rect 273694 82294 273762 82350
rect 273818 82294 273888 82350
rect 273568 82226 273888 82294
rect 273568 82170 273638 82226
rect 273694 82170 273762 82226
rect 273818 82170 273888 82226
rect 273568 82102 273888 82170
rect 273568 82046 273638 82102
rect 273694 82046 273762 82102
rect 273818 82046 273888 82102
rect 273568 81978 273888 82046
rect 273568 81922 273638 81978
rect 273694 81922 273762 81978
rect 273818 81922 273888 81978
rect 273568 81888 273888 81922
rect 304288 82350 304608 82384
rect 304288 82294 304358 82350
rect 304414 82294 304482 82350
rect 304538 82294 304608 82350
rect 304288 82226 304608 82294
rect 304288 82170 304358 82226
rect 304414 82170 304482 82226
rect 304538 82170 304608 82226
rect 304288 82102 304608 82170
rect 304288 82046 304358 82102
rect 304414 82046 304482 82102
rect 304538 82046 304608 82102
rect 304288 81978 304608 82046
rect 304288 81922 304358 81978
rect 304414 81922 304482 81978
rect 304538 81922 304608 81978
rect 304288 81888 304608 81922
rect 335008 82350 335328 82384
rect 335008 82294 335078 82350
rect 335134 82294 335202 82350
rect 335258 82294 335328 82350
rect 335008 82226 335328 82294
rect 335008 82170 335078 82226
rect 335134 82170 335202 82226
rect 335258 82170 335328 82226
rect 335008 82102 335328 82170
rect 335008 82046 335078 82102
rect 335134 82046 335202 82102
rect 335258 82046 335328 82102
rect 335008 81978 335328 82046
rect 335008 81922 335078 81978
rect 335134 81922 335202 81978
rect 335258 81922 335328 81978
rect 335008 81888 335328 81922
rect 365728 82350 366048 82384
rect 365728 82294 365798 82350
rect 365854 82294 365922 82350
rect 365978 82294 366048 82350
rect 365728 82226 366048 82294
rect 365728 82170 365798 82226
rect 365854 82170 365922 82226
rect 365978 82170 366048 82226
rect 365728 82102 366048 82170
rect 365728 82046 365798 82102
rect 365854 82046 365922 82102
rect 365978 82046 366048 82102
rect 365728 81978 366048 82046
rect 365728 81922 365798 81978
rect 365854 81922 365922 81978
rect 365978 81922 366048 81978
rect 365728 81888 366048 81922
rect 396448 82350 396768 82384
rect 396448 82294 396518 82350
rect 396574 82294 396642 82350
rect 396698 82294 396768 82350
rect 396448 82226 396768 82294
rect 396448 82170 396518 82226
rect 396574 82170 396642 82226
rect 396698 82170 396768 82226
rect 396448 82102 396768 82170
rect 396448 82046 396518 82102
rect 396574 82046 396642 82102
rect 396698 82046 396768 82102
rect 396448 81978 396768 82046
rect 396448 81922 396518 81978
rect 396574 81922 396642 81978
rect 396698 81922 396768 81978
rect 396448 81888 396768 81922
rect 427168 82350 427488 82384
rect 427168 82294 427238 82350
rect 427294 82294 427362 82350
rect 427418 82294 427488 82350
rect 427168 82226 427488 82294
rect 427168 82170 427238 82226
rect 427294 82170 427362 82226
rect 427418 82170 427488 82226
rect 427168 82102 427488 82170
rect 427168 82046 427238 82102
rect 427294 82046 427362 82102
rect 427418 82046 427488 82102
rect 427168 81978 427488 82046
rect 427168 81922 427238 81978
rect 427294 81922 427362 81978
rect 427418 81922 427488 81978
rect 427168 81888 427488 81922
rect 457888 82350 458208 82384
rect 457888 82294 457958 82350
rect 458014 82294 458082 82350
rect 458138 82294 458208 82350
rect 457888 82226 458208 82294
rect 457888 82170 457958 82226
rect 458014 82170 458082 82226
rect 458138 82170 458208 82226
rect 457888 82102 458208 82170
rect 457888 82046 457958 82102
rect 458014 82046 458082 82102
rect 458138 82046 458208 82102
rect 457888 81978 458208 82046
rect 457888 81922 457958 81978
rect 458014 81922 458082 81978
rect 458138 81922 458208 81978
rect 457888 81888 458208 81922
rect 488608 82350 488928 82384
rect 488608 82294 488678 82350
rect 488734 82294 488802 82350
rect 488858 82294 488928 82350
rect 488608 82226 488928 82294
rect 488608 82170 488678 82226
rect 488734 82170 488802 82226
rect 488858 82170 488928 82226
rect 488608 82102 488928 82170
rect 488608 82046 488678 82102
rect 488734 82046 488802 82102
rect 488858 82046 488928 82102
rect 488608 81978 488928 82046
rect 488608 81922 488678 81978
rect 488734 81922 488802 81978
rect 488858 81922 488928 81978
rect 488608 81888 488928 81922
rect 519328 82350 519648 82384
rect 519328 82294 519398 82350
rect 519454 82294 519522 82350
rect 519578 82294 519648 82350
rect 519328 82226 519648 82294
rect 519328 82170 519398 82226
rect 519454 82170 519522 82226
rect 519578 82170 519648 82226
rect 519328 82102 519648 82170
rect 519328 82046 519398 82102
rect 519454 82046 519522 82102
rect 519578 82046 519648 82102
rect 519328 81978 519648 82046
rect 519328 81922 519398 81978
rect 519454 81922 519522 81978
rect 519578 81922 519648 81978
rect 519328 81888 519648 81922
rect 550048 82350 550368 82384
rect 550048 82294 550118 82350
rect 550174 82294 550242 82350
rect 550298 82294 550368 82350
rect 550048 82226 550368 82294
rect 550048 82170 550118 82226
rect 550174 82170 550242 82226
rect 550298 82170 550368 82226
rect 550048 82102 550368 82170
rect 550048 82046 550118 82102
rect 550174 82046 550242 82102
rect 550298 82046 550368 82102
rect 550048 81978 550368 82046
rect 550048 81922 550118 81978
rect 550174 81922 550242 81978
rect 550298 81922 550368 81978
rect 550048 81888 550368 81922
rect 5418 76294 5514 76350
rect 5570 76294 5638 76350
rect 5694 76294 5762 76350
rect 5818 76294 5886 76350
rect 5942 76294 6038 76350
rect 5418 76226 6038 76294
rect 5418 76170 5514 76226
rect 5570 76170 5638 76226
rect 5694 76170 5762 76226
rect 5818 76170 5886 76226
rect 5942 76170 6038 76226
rect 5418 76102 6038 76170
rect 5418 76046 5514 76102
rect 5570 76046 5638 76102
rect 5694 76046 5762 76102
rect 5818 76046 5886 76102
rect 5942 76046 6038 76102
rect 5418 75978 6038 76046
rect 5418 75922 5514 75978
rect 5570 75922 5638 75978
rect 5694 75922 5762 75978
rect 5818 75922 5886 75978
rect 5942 75922 6038 75978
rect 5068 65044 5124 65054
rect 5068 59780 5124 64988
rect 5068 59714 5124 59724
rect -956 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 -336 58350
rect -956 58226 -336 58294
rect -956 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 -336 58226
rect -956 58102 -336 58170
rect -956 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 -336 58102
rect -956 57978 -336 58046
rect -956 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 -336 57978
rect -956 40350 -336 57922
rect 5418 58350 6038 75922
rect 12448 76350 12768 76384
rect 12448 76294 12518 76350
rect 12574 76294 12642 76350
rect 12698 76294 12768 76350
rect 12448 76226 12768 76294
rect 12448 76170 12518 76226
rect 12574 76170 12642 76226
rect 12698 76170 12768 76226
rect 12448 76102 12768 76170
rect 12448 76046 12518 76102
rect 12574 76046 12642 76102
rect 12698 76046 12768 76102
rect 12448 75978 12768 76046
rect 12448 75922 12518 75978
rect 12574 75922 12642 75978
rect 12698 75922 12768 75978
rect 12448 75888 12768 75922
rect 43168 76350 43488 76384
rect 43168 76294 43238 76350
rect 43294 76294 43362 76350
rect 43418 76294 43488 76350
rect 43168 76226 43488 76294
rect 43168 76170 43238 76226
rect 43294 76170 43362 76226
rect 43418 76170 43488 76226
rect 43168 76102 43488 76170
rect 43168 76046 43238 76102
rect 43294 76046 43362 76102
rect 43418 76046 43488 76102
rect 43168 75978 43488 76046
rect 43168 75922 43238 75978
rect 43294 75922 43362 75978
rect 43418 75922 43488 75978
rect 43168 75888 43488 75922
rect 73888 76350 74208 76384
rect 73888 76294 73958 76350
rect 74014 76294 74082 76350
rect 74138 76294 74208 76350
rect 73888 76226 74208 76294
rect 73888 76170 73958 76226
rect 74014 76170 74082 76226
rect 74138 76170 74208 76226
rect 73888 76102 74208 76170
rect 73888 76046 73958 76102
rect 74014 76046 74082 76102
rect 74138 76046 74208 76102
rect 73888 75978 74208 76046
rect 73888 75922 73958 75978
rect 74014 75922 74082 75978
rect 74138 75922 74208 75978
rect 73888 75888 74208 75922
rect 104608 76350 104928 76384
rect 104608 76294 104678 76350
rect 104734 76294 104802 76350
rect 104858 76294 104928 76350
rect 104608 76226 104928 76294
rect 104608 76170 104678 76226
rect 104734 76170 104802 76226
rect 104858 76170 104928 76226
rect 104608 76102 104928 76170
rect 104608 76046 104678 76102
rect 104734 76046 104802 76102
rect 104858 76046 104928 76102
rect 104608 75978 104928 76046
rect 104608 75922 104678 75978
rect 104734 75922 104802 75978
rect 104858 75922 104928 75978
rect 104608 75888 104928 75922
rect 135328 76350 135648 76384
rect 135328 76294 135398 76350
rect 135454 76294 135522 76350
rect 135578 76294 135648 76350
rect 135328 76226 135648 76294
rect 135328 76170 135398 76226
rect 135454 76170 135522 76226
rect 135578 76170 135648 76226
rect 135328 76102 135648 76170
rect 135328 76046 135398 76102
rect 135454 76046 135522 76102
rect 135578 76046 135648 76102
rect 135328 75978 135648 76046
rect 135328 75922 135398 75978
rect 135454 75922 135522 75978
rect 135578 75922 135648 75978
rect 135328 75888 135648 75922
rect 166048 76350 166368 76384
rect 166048 76294 166118 76350
rect 166174 76294 166242 76350
rect 166298 76294 166368 76350
rect 166048 76226 166368 76294
rect 166048 76170 166118 76226
rect 166174 76170 166242 76226
rect 166298 76170 166368 76226
rect 166048 76102 166368 76170
rect 166048 76046 166118 76102
rect 166174 76046 166242 76102
rect 166298 76046 166368 76102
rect 166048 75978 166368 76046
rect 166048 75922 166118 75978
rect 166174 75922 166242 75978
rect 166298 75922 166368 75978
rect 166048 75888 166368 75922
rect 196768 76350 197088 76384
rect 196768 76294 196838 76350
rect 196894 76294 196962 76350
rect 197018 76294 197088 76350
rect 196768 76226 197088 76294
rect 196768 76170 196838 76226
rect 196894 76170 196962 76226
rect 197018 76170 197088 76226
rect 196768 76102 197088 76170
rect 196768 76046 196838 76102
rect 196894 76046 196962 76102
rect 197018 76046 197088 76102
rect 196768 75978 197088 76046
rect 196768 75922 196838 75978
rect 196894 75922 196962 75978
rect 197018 75922 197088 75978
rect 196768 75888 197088 75922
rect 227488 76350 227808 76384
rect 227488 76294 227558 76350
rect 227614 76294 227682 76350
rect 227738 76294 227808 76350
rect 227488 76226 227808 76294
rect 227488 76170 227558 76226
rect 227614 76170 227682 76226
rect 227738 76170 227808 76226
rect 227488 76102 227808 76170
rect 227488 76046 227558 76102
rect 227614 76046 227682 76102
rect 227738 76046 227808 76102
rect 227488 75978 227808 76046
rect 227488 75922 227558 75978
rect 227614 75922 227682 75978
rect 227738 75922 227808 75978
rect 227488 75888 227808 75922
rect 258208 76350 258528 76384
rect 258208 76294 258278 76350
rect 258334 76294 258402 76350
rect 258458 76294 258528 76350
rect 258208 76226 258528 76294
rect 258208 76170 258278 76226
rect 258334 76170 258402 76226
rect 258458 76170 258528 76226
rect 258208 76102 258528 76170
rect 258208 76046 258278 76102
rect 258334 76046 258402 76102
rect 258458 76046 258528 76102
rect 258208 75978 258528 76046
rect 258208 75922 258278 75978
rect 258334 75922 258402 75978
rect 258458 75922 258528 75978
rect 258208 75888 258528 75922
rect 288928 76350 289248 76384
rect 288928 76294 288998 76350
rect 289054 76294 289122 76350
rect 289178 76294 289248 76350
rect 288928 76226 289248 76294
rect 288928 76170 288998 76226
rect 289054 76170 289122 76226
rect 289178 76170 289248 76226
rect 288928 76102 289248 76170
rect 288928 76046 288998 76102
rect 289054 76046 289122 76102
rect 289178 76046 289248 76102
rect 288928 75978 289248 76046
rect 288928 75922 288998 75978
rect 289054 75922 289122 75978
rect 289178 75922 289248 75978
rect 288928 75888 289248 75922
rect 319648 76350 319968 76384
rect 319648 76294 319718 76350
rect 319774 76294 319842 76350
rect 319898 76294 319968 76350
rect 319648 76226 319968 76294
rect 319648 76170 319718 76226
rect 319774 76170 319842 76226
rect 319898 76170 319968 76226
rect 319648 76102 319968 76170
rect 319648 76046 319718 76102
rect 319774 76046 319842 76102
rect 319898 76046 319968 76102
rect 319648 75978 319968 76046
rect 319648 75922 319718 75978
rect 319774 75922 319842 75978
rect 319898 75922 319968 75978
rect 319648 75888 319968 75922
rect 350368 76350 350688 76384
rect 350368 76294 350438 76350
rect 350494 76294 350562 76350
rect 350618 76294 350688 76350
rect 350368 76226 350688 76294
rect 350368 76170 350438 76226
rect 350494 76170 350562 76226
rect 350618 76170 350688 76226
rect 350368 76102 350688 76170
rect 350368 76046 350438 76102
rect 350494 76046 350562 76102
rect 350618 76046 350688 76102
rect 350368 75978 350688 76046
rect 350368 75922 350438 75978
rect 350494 75922 350562 75978
rect 350618 75922 350688 75978
rect 350368 75888 350688 75922
rect 381088 76350 381408 76384
rect 381088 76294 381158 76350
rect 381214 76294 381282 76350
rect 381338 76294 381408 76350
rect 381088 76226 381408 76294
rect 381088 76170 381158 76226
rect 381214 76170 381282 76226
rect 381338 76170 381408 76226
rect 381088 76102 381408 76170
rect 381088 76046 381158 76102
rect 381214 76046 381282 76102
rect 381338 76046 381408 76102
rect 381088 75978 381408 76046
rect 381088 75922 381158 75978
rect 381214 75922 381282 75978
rect 381338 75922 381408 75978
rect 381088 75888 381408 75922
rect 411808 76350 412128 76384
rect 411808 76294 411878 76350
rect 411934 76294 412002 76350
rect 412058 76294 412128 76350
rect 411808 76226 412128 76294
rect 411808 76170 411878 76226
rect 411934 76170 412002 76226
rect 412058 76170 412128 76226
rect 411808 76102 412128 76170
rect 411808 76046 411878 76102
rect 411934 76046 412002 76102
rect 412058 76046 412128 76102
rect 411808 75978 412128 76046
rect 411808 75922 411878 75978
rect 411934 75922 412002 75978
rect 412058 75922 412128 75978
rect 411808 75888 412128 75922
rect 442528 76350 442848 76384
rect 442528 76294 442598 76350
rect 442654 76294 442722 76350
rect 442778 76294 442848 76350
rect 442528 76226 442848 76294
rect 442528 76170 442598 76226
rect 442654 76170 442722 76226
rect 442778 76170 442848 76226
rect 442528 76102 442848 76170
rect 442528 76046 442598 76102
rect 442654 76046 442722 76102
rect 442778 76046 442848 76102
rect 442528 75978 442848 76046
rect 442528 75922 442598 75978
rect 442654 75922 442722 75978
rect 442778 75922 442848 75978
rect 442528 75888 442848 75922
rect 473248 76350 473568 76384
rect 473248 76294 473318 76350
rect 473374 76294 473442 76350
rect 473498 76294 473568 76350
rect 473248 76226 473568 76294
rect 473248 76170 473318 76226
rect 473374 76170 473442 76226
rect 473498 76170 473568 76226
rect 473248 76102 473568 76170
rect 473248 76046 473318 76102
rect 473374 76046 473442 76102
rect 473498 76046 473568 76102
rect 473248 75978 473568 76046
rect 473248 75922 473318 75978
rect 473374 75922 473442 75978
rect 473498 75922 473568 75978
rect 473248 75888 473568 75922
rect 503968 76350 504288 76384
rect 503968 76294 504038 76350
rect 504094 76294 504162 76350
rect 504218 76294 504288 76350
rect 503968 76226 504288 76294
rect 503968 76170 504038 76226
rect 504094 76170 504162 76226
rect 504218 76170 504288 76226
rect 503968 76102 504288 76170
rect 503968 76046 504038 76102
rect 504094 76046 504162 76102
rect 504218 76046 504288 76102
rect 503968 75978 504288 76046
rect 503968 75922 504038 75978
rect 504094 75922 504162 75978
rect 504218 75922 504288 75978
rect 503968 75888 504288 75922
rect 534688 76350 535008 76384
rect 534688 76294 534758 76350
rect 534814 76294 534882 76350
rect 534938 76294 535008 76350
rect 534688 76226 535008 76294
rect 534688 76170 534758 76226
rect 534814 76170 534882 76226
rect 534938 76170 535008 76226
rect 534688 76102 535008 76170
rect 534688 76046 534758 76102
rect 534814 76046 534882 76102
rect 534938 76046 535008 76102
rect 534688 75978 535008 76046
rect 534688 75922 534758 75978
rect 534814 75922 534882 75978
rect 534938 75922 535008 75978
rect 534688 75888 535008 75922
rect 565408 76350 565728 76384
rect 565408 76294 565478 76350
rect 565534 76294 565602 76350
rect 565658 76294 565728 76350
rect 565408 76226 565728 76294
rect 565408 76170 565478 76226
rect 565534 76170 565602 76226
rect 565658 76170 565728 76226
rect 565408 76102 565728 76170
rect 565408 76046 565478 76102
rect 565534 76046 565602 76102
rect 565658 76046 565728 76102
rect 565408 75978 565728 76046
rect 565408 75922 565478 75978
rect 565534 75922 565602 75978
rect 565658 75922 565728 75978
rect 565408 75888 565728 75922
rect 589098 76350 589718 93922
rect 592818 100350 593438 117922
rect 592818 100294 592914 100350
rect 592970 100294 593038 100350
rect 593094 100294 593162 100350
rect 593218 100294 593286 100350
rect 593342 100294 593438 100350
rect 592818 100226 593438 100294
rect 592818 100170 592914 100226
rect 592970 100170 593038 100226
rect 593094 100170 593162 100226
rect 593218 100170 593286 100226
rect 593342 100170 593438 100226
rect 592818 100102 593438 100170
rect 592818 100046 592914 100102
rect 592970 100046 593038 100102
rect 593094 100046 593162 100102
rect 593218 100046 593286 100102
rect 593342 100046 593438 100102
rect 592818 99978 593438 100046
rect 592818 99922 592914 99978
rect 592970 99922 593038 99978
rect 593094 99922 593162 99978
rect 593218 99922 593286 99978
rect 593342 99922 593438 99978
rect 590492 86436 590548 86446
rect 590492 81732 590548 86380
rect 590492 81666 590548 81676
rect 592818 82350 593438 99922
rect 592818 82294 592914 82350
rect 592970 82294 593038 82350
rect 593094 82294 593162 82350
rect 593218 82294 593286 82350
rect 593342 82294 593438 82350
rect 592818 82226 593438 82294
rect 592818 82170 592914 82226
rect 592970 82170 593038 82226
rect 593094 82170 593162 82226
rect 593218 82170 593286 82226
rect 593342 82170 593438 82226
rect 592818 82102 593438 82170
rect 592818 82046 592914 82102
rect 592970 82046 593038 82102
rect 593094 82046 593162 82102
rect 593218 82046 593286 82102
rect 593342 82046 593438 82102
rect 592818 81978 593438 82046
rect 592818 81922 592914 81978
rect 592970 81922 593038 81978
rect 593094 81922 593162 81978
rect 593218 81922 593286 81978
rect 593342 81922 593438 81978
rect 589098 76294 589194 76350
rect 589250 76294 589318 76350
rect 589374 76294 589442 76350
rect 589498 76294 589566 76350
rect 589622 76294 589718 76350
rect 589098 76226 589718 76294
rect 589098 76170 589194 76226
rect 589250 76170 589318 76226
rect 589374 76170 589442 76226
rect 589498 76170 589566 76226
rect 589622 76170 589718 76226
rect 589098 76102 589718 76170
rect 589098 76046 589194 76102
rect 589250 76046 589318 76102
rect 589374 76046 589442 76102
rect 589498 76046 589566 76102
rect 589622 76046 589718 76102
rect 589098 75978 589718 76046
rect 589098 75922 589194 75978
rect 589250 75922 589318 75978
rect 589374 75922 589442 75978
rect 589498 75922 589566 75978
rect 589622 75922 589718 75978
rect 588924 73220 588980 73230
rect 588924 70980 588980 73164
rect 588924 70914 588980 70924
rect 27808 64350 28128 64384
rect 27808 64294 27878 64350
rect 27934 64294 28002 64350
rect 28058 64294 28128 64350
rect 27808 64226 28128 64294
rect 27808 64170 27878 64226
rect 27934 64170 28002 64226
rect 28058 64170 28128 64226
rect 27808 64102 28128 64170
rect 27808 64046 27878 64102
rect 27934 64046 28002 64102
rect 28058 64046 28128 64102
rect 27808 63978 28128 64046
rect 27808 63922 27878 63978
rect 27934 63922 28002 63978
rect 28058 63922 28128 63978
rect 27808 63888 28128 63922
rect 58528 64350 58848 64384
rect 58528 64294 58598 64350
rect 58654 64294 58722 64350
rect 58778 64294 58848 64350
rect 58528 64226 58848 64294
rect 58528 64170 58598 64226
rect 58654 64170 58722 64226
rect 58778 64170 58848 64226
rect 58528 64102 58848 64170
rect 58528 64046 58598 64102
rect 58654 64046 58722 64102
rect 58778 64046 58848 64102
rect 58528 63978 58848 64046
rect 58528 63922 58598 63978
rect 58654 63922 58722 63978
rect 58778 63922 58848 63978
rect 58528 63888 58848 63922
rect 89248 64350 89568 64384
rect 89248 64294 89318 64350
rect 89374 64294 89442 64350
rect 89498 64294 89568 64350
rect 89248 64226 89568 64294
rect 89248 64170 89318 64226
rect 89374 64170 89442 64226
rect 89498 64170 89568 64226
rect 89248 64102 89568 64170
rect 89248 64046 89318 64102
rect 89374 64046 89442 64102
rect 89498 64046 89568 64102
rect 89248 63978 89568 64046
rect 89248 63922 89318 63978
rect 89374 63922 89442 63978
rect 89498 63922 89568 63978
rect 89248 63888 89568 63922
rect 119968 64350 120288 64384
rect 119968 64294 120038 64350
rect 120094 64294 120162 64350
rect 120218 64294 120288 64350
rect 119968 64226 120288 64294
rect 119968 64170 120038 64226
rect 120094 64170 120162 64226
rect 120218 64170 120288 64226
rect 119968 64102 120288 64170
rect 119968 64046 120038 64102
rect 120094 64046 120162 64102
rect 120218 64046 120288 64102
rect 119968 63978 120288 64046
rect 119968 63922 120038 63978
rect 120094 63922 120162 63978
rect 120218 63922 120288 63978
rect 119968 63888 120288 63922
rect 150688 64350 151008 64384
rect 150688 64294 150758 64350
rect 150814 64294 150882 64350
rect 150938 64294 151008 64350
rect 150688 64226 151008 64294
rect 150688 64170 150758 64226
rect 150814 64170 150882 64226
rect 150938 64170 151008 64226
rect 150688 64102 151008 64170
rect 150688 64046 150758 64102
rect 150814 64046 150882 64102
rect 150938 64046 151008 64102
rect 150688 63978 151008 64046
rect 150688 63922 150758 63978
rect 150814 63922 150882 63978
rect 150938 63922 151008 63978
rect 150688 63888 151008 63922
rect 181408 64350 181728 64384
rect 181408 64294 181478 64350
rect 181534 64294 181602 64350
rect 181658 64294 181728 64350
rect 181408 64226 181728 64294
rect 181408 64170 181478 64226
rect 181534 64170 181602 64226
rect 181658 64170 181728 64226
rect 181408 64102 181728 64170
rect 181408 64046 181478 64102
rect 181534 64046 181602 64102
rect 181658 64046 181728 64102
rect 181408 63978 181728 64046
rect 181408 63922 181478 63978
rect 181534 63922 181602 63978
rect 181658 63922 181728 63978
rect 181408 63888 181728 63922
rect 212128 64350 212448 64384
rect 212128 64294 212198 64350
rect 212254 64294 212322 64350
rect 212378 64294 212448 64350
rect 212128 64226 212448 64294
rect 212128 64170 212198 64226
rect 212254 64170 212322 64226
rect 212378 64170 212448 64226
rect 212128 64102 212448 64170
rect 212128 64046 212198 64102
rect 212254 64046 212322 64102
rect 212378 64046 212448 64102
rect 212128 63978 212448 64046
rect 212128 63922 212198 63978
rect 212254 63922 212322 63978
rect 212378 63922 212448 63978
rect 212128 63888 212448 63922
rect 242848 64350 243168 64384
rect 242848 64294 242918 64350
rect 242974 64294 243042 64350
rect 243098 64294 243168 64350
rect 242848 64226 243168 64294
rect 242848 64170 242918 64226
rect 242974 64170 243042 64226
rect 243098 64170 243168 64226
rect 242848 64102 243168 64170
rect 242848 64046 242918 64102
rect 242974 64046 243042 64102
rect 243098 64046 243168 64102
rect 242848 63978 243168 64046
rect 242848 63922 242918 63978
rect 242974 63922 243042 63978
rect 243098 63922 243168 63978
rect 242848 63888 243168 63922
rect 273568 64350 273888 64384
rect 273568 64294 273638 64350
rect 273694 64294 273762 64350
rect 273818 64294 273888 64350
rect 273568 64226 273888 64294
rect 273568 64170 273638 64226
rect 273694 64170 273762 64226
rect 273818 64170 273888 64226
rect 273568 64102 273888 64170
rect 273568 64046 273638 64102
rect 273694 64046 273762 64102
rect 273818 64046 273888 64102
rect 273568 63978 273888 64046
rect 273568 63922 273638 63978
rect 273694 63922 273762 63978
rect 273818 63922 273888 63978
rect 273568 63888 273888 63922
rect 304288 64350 304608 64384
rect 304288 64294 304358 64350
rect 304414 64294 304482 64350
rect 304538 64294 304608 64350
rect 304288 64226 304608 64294
rect 304288 64170 304358 64226
rect 304414 64170 304482 64226
rect 304538 64170 304608 64226
rect 304288 64102 304608 64170
rect 304288 64046 304358 64102
rect 304414 64046 304482 64102
rect 304538 64046 304608 64102
rect 304288 63978 304608 64046
rect 304288 63922 304358 63978
rect 304414 63922 304482 63978
rect 304538 63922 304608 63978
rect 304288 63888 304608 63922
rect 335008 64350 335328 64384
rect 335008 64294 335078 64350
rect 335134 64294 335202 64350
rect 335258 64294 335328 64350
rect 335008 64226 335328 64294
rect 335008 64170 335078 64226
rect 335134 64170 335202 64226
rect 335258 64170 335328 64226
rect 335008 64102 335328 64170
rect 335008 64046 335078 64102
rect 335134 64046 335202 64102
rect 335258 64046 335328 64102
rect 335008 63978 335328 64046
rect 335008 63922 335078 63978
rect 335134 63922 335202 63978
rect 335258 63922 335328 63978
rect 335008 63888 335328 63922
rect 365728 64350 366048 64384
rect 365728 64294 365798 64350
rect 365854 64294 365922 64350
rect 365978 64294 366048 64350
rect 365728 64226 366048 64294
rect 365728 64170 365798 64226
rect 365854 64170 365922 64226
rect 365978 64170 366048 64226
rect 365728 64102 366048 64170
rect 365728 64046 365798 64102
rect 365854 64046 365922 64102
rect 365978 64046 366048 64102
rect 365728 63978 366048 64046
rect 365728 63922 365798 63978
rect 365854 63922 365922 63978
rect 365978 63922 366048 63978
rect 365728 63888 366048 63922
rect 396448 64350 396768 64384
rect 396448 64294 396518 64350
rect 396574 64294 396642 64350
rect 396698 64294 396768 64350
rect 396448 64226 396768 64294
rect 396448 64170 396518 64226
rect 396574 64170 396642 64226
rect 396698 64170 396768 64226
rect 396448 64102 396768 64170
rect 396448 64046 396518 64102
rect 396574 64046 396642 64102
rect 396698 64046 396768 64102
rect 396448 63978 396768 64046
rect 396448 63922 396518 63978
rect 396574 63922 396642 63978
rect 396698 63922 396768 63978
rect 396448 63888 396768 63922
rect 427168 64350 427488 64384
rect 427168 64294 427238 64350
rect 427294 64294 427362 64350
rect 427418 64294 427488 64350
rect 427168 64226 427488 64294
rect 427168 64170 427238 64226
rect 427294 64170 427362 64226
rect 427418 64170 427488 64226
rect 427168 64102 427488 64170
rect 427168 64046 427238 64102
rect 427294 64046 427362 64102
rect 427418 64046 427488 64102
rect 427168 63978 427488 64046
rect 427168 63922 427238 63978
rect 427294 63922 427362 63978
rect 427418 63922 427488 63978
rect 427168 63888 427488 63922
rect 457888 64350 458208 64384
rect 457888 64294 457958 64350
rect 458014 64294 458082 64350
rect 458138 64294 458208 64350
rect 457888 64226 458208 64294
rect 457888 64170 457958 64226
rect 458014 64170 458082 64226
rect 458138 64170 458208 64226
rect 457888 64102 458208 64170
rect 457888 64046 457958 64102
rect 458014 64046 458082 64102
rect 458138 64046 458208 64102
rect 457888 63978 458208 64046
rect 457888 63922 457958 63978
rect 458014 63922 458082 63978
rect 458138 63922 458208 63978
rect 457888 63888 458208 63922
rect 488608 64350 488928 64384
rect 488608 64294 488678 64350
rect 488734 64294 488802 64350
rect 488858 64294 488928 64350
rect 488608 64226 488928 64294
rect 488608 64170 488678 64226
rect 488734 64170 488802 64226
rect 488858 64170 488928 64226
rect 488608 64102 488928 64170
rect 488608 64046 488678 64102
rect 488734 64046 488802 64102
rect 488858 64046 488928 64102
rect 488608 63978 488928 64046
rect 488608 63922 488678 63978
rect 488734 63922 488802 63978
rect 488858 63922 488928 63978
rect 488608 63888 488928 63922
rect 519328 64350 519648 64384
rect 519328 64294 519398 64350
rect 519454 64294 519522 64350
rect 519578 64294 519648 64350
rect 519328 64226 519648 64294
rect 519328 64170 519398 64226
rect 519454 64170 519522 64226
rect 519578 64170 519648 64226
rect 519328 64102 519648 64170
rect 519328 64046 519398 64102
rect 519454 64046 519522 64102
rect 519578 64046 519648 64102
rect 519328 63978 519648 64046
rect 519328 63922 519398 63978
rect 519454 63922 519522 63978
rect 519578 63922 519648 63978
rect 519328 63888 519648 63922
rect 550048 64350 550368 64384
rect 550048 64294 550118 64350
rect 550174 64294 550242 64350
rect 550298 64294 550368 64350
rect 550048 64226 550368 64294
rect 550048 64170 550118 64226
rect 550174 64170 550242 64226
rect 550298 64170 550368 64226
rect 550048 64102 550368 64170
rect 550048 64046 550118 64102
rect 550174 64046 550242 64102
rect 550298 64046 550368 64102
rect 550048 63978 550368 64046
rect 550048 63922 550118 63978
rect 550174 63922 550242 63978
rect 550298 63922 550368 63978
rect 550048 63888 550368 63922
rect 5418 58294 5514 58350
rect 5570 58294 5638 58350
rect 5694 58294 5762 58350
rect 5818 58294 5886 58350
rect 5942 58294 6038 58350
rect 5418 58226 6038 58294
rect 5418 58170 5514 58226
rect 5570 58170 5638 58226
rect 5694 58170 5762 58226
rect 5818 58170 5886 58226
rect 5942 58170 6038 58226
rect 5418 58102 6038 58170
rect 5418 58046 5514 58102
rect 5570 58046 5638 58102
rect 5694 58046 5762 58102
rect 5818 58046 5886 58102
rect 5942 58046 6038 58102
rect 5418 57978 6038 58046
rect 5418 57922 5514 57978
rect 5570 57922 5638 57978
rect 5694 57922 5762 57978
rect 5818 57922 5886 57978
rect 5942 57922 6038 57978
rect 5068 50932 5124 50942
rect 5068 49252 5124 50876
rect 5068 49186 5124 49196
rect -956 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 -336 40350
rect -956 40226 -336 40294
rect -956 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 -336 40226
rect -956 40102 -336 40170
rect -956 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 -336 40102
rect -956 39978 -336 40046
rect -956 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 -336 39978
rect -956 22350 -336 39922
rect 5418 40350 6038 57922
rect 12448 58350 12768 58384
rect 12448 58294 12518 58350
rect 12574 58294 12642 58350
rect 12698 58294 12768 58350
rect 12448 58226 12768 58294
rect 12448 58170 12518 58226
rect 12574 58170 12642 58226
rect 12698 58170 12768 58226
rect 12448 58102 12768 58170
rect 12448 58046 12518 58102
rect 12574 58046 12642 58102
rect 12698 58046 12768 58102
rect 12448 57978 12768 58046
rect 12448 57922 12518 57978
rect 12574 57922 12642 57978
rect 12698 57922 12768 57978
rect 12448 57888 12768 57922
rect 43168 58350 43488 58384
rect 43168 58294 43238 58350
rect 43294 58294 43362 58350
rect 43418 58294 43488 58350
rect 43168 58226 43488 58294
rect 43168 58170 43238 58226
rect 43294 58170 43362 58226
rect 43418 58170 43488 58226
rect 43168 58102 43488 58170
rect 43168 58046 43238 58102
rect 43294 58046 43362 58102
rect 43418 58046 43488 58102
rect 43168 57978 43488 58046
rect 43168 57922 43238 57978
rect 43294 57922 43362 57978
rect 43418 57922 43488 57978
rect 43168 57888 43488 57922
rect 73888 58350 74208 58384
rect 73888 58294 73958 58350
rect 74014 58294 74082 58350
rect 74138 58294 74208 58350
rect 73888 58226 74208 58294
rect 73888 58170 73958 58226
rect 74014 58170 74082 58226
rect 74138 58170 74208 58226
rect 73888 58102 74208 58170
rect 73888 58046 73958 58102
rect 74014 58046 74082 58102
rect 74138 58046 74208 58102
rect 73888 57978 74208 58046
rect 73888 57922 73958 57978
rect 74014 57922 74082 57978
rect 74138 57922 74208 57978
rect 73888 57888 74208 57922
rect 104608 58350 104928 58384
rect 104608 58294 104678 58350
rect 104734 58294 104802 58350
rect 104858 58294 104928 58350
rect 104608 58226 104928 58294
rect 104608 58170 104678 58226
rect 104734 58170 104802 58226
rect 104858 58170 104928 58226
rect 104608 58102 104928 58170
rect 104608 58046 104678 58102
rect 104734 58046 104802 58102
rect 104858 58046 104928 58102
rect 104608 57978 104928 58046
rect 104608 57922 104678 57978
rect 104734 57922 104802 57978
rect 104858 57922 104928 57978
rect 104608 57888 104928 57922
rect 135328 58350 135648 58384
rect 135328 58294 135398 58350
rect 135454 58294 135522 58350
rect 135578 58294 135648 58350
rect 135328 58226 135648 58294
rect 135328 58170 135398 58226
rect 135454 58170 135522 58226
rect 135578 58170 135648 58226
rect 135328 58102 135648 58170
rect 135328 58046 135398 58102
rect 135454 58046 135522 58102
rect 135578 58046 135648 58102
rect 135328 57978 135648 58046
rect 135328 57922 135398 57978
rect 135454 57922 135522 57978
rect 135578 57922 135648 57978
rect 135328 57888 135648 57922
rect 166048 58350 166368 58384
rect 166048 58294 166118 58350
rect 166174 58294 166242 58350
rect 166298 58294 166368 58350
rect 166048 58226 166368 58294
rect 166048 58170 166118 58226
rect 166174 58170 166242 58226
rect 166298 58170 166368 58226
rect 166048 58102 166368 58170
rect 166048 58046 166118 58102
rect 166174 58046 166242 58102
rect 166298 58046 166368 58102
rect 166048 57978 166368 58046
rect 166048 57922 166118 57978
rect 166174 57922 166242 57978
rect 166298 57922 166368 57978
rect 166048 57888 166368 57922
rect 196768 58350 197088 58384
rect 196768 58294 196838 58350
rect 196894 58294 196962 58350
rect 197018 58294 197088 58350
rect 196768 58226 197088 58294
rect 196768 58170 196838 58226
rect 196894 58170 196962 58226
rect 197018 58170 197088 58226
rect 196768 58102 197088 58170
rect 196768 58046 196838 58102
rect 196894 58046 196962 58102
rect 197018 58046 197088 58102
rect 196768 57978 197088 58046
rect 196768 57922 196838 57978
rect 196894 57922 196962 57978
rect 197018 57922 197088 57978
rect 196768 57888 197088 57922
rect 227488 58350 227808 58384
rect 227488 58294 227558 58350
rect 227614 58294 227682 58350
rect 227738 58294 227808 58350
rect 227488 58226 227808 58294
rect 227488 58170 227558 58226
rect 227614 58170 227682 58226
rect 227738 58170 227808 58226
rect 227488 58102 227808 58170
rect 227488 58046 227558 58102
rect 227614 58046 227682 58102
rect 227738 58046 227808 58102
rect 227488 57978 227808 58046
rect 227488 57922 227558 57978
rect 227614 57922 227682 57978
rect 227738 57922 227808 57978
rect 227488 57888 227808 57922
rect 258208 58350 258528 58384
rect 258208 58294 258278 58350
rect 258334 58294 258402 58350
rect 258458 58294 258528 58350
rect 258208 58226 258528 58294
rect 258208 58170 258278 58226
rect 258334 58170 258402 58226
rect 258458 58170 258528 58226
rect 258208 58102 258528 58170
rect 258208 58046 258278 58102
rect 258334 58046 258402 58102
rect 258458 58046 258528 58102
rect 258208 57978 258528 58046
rect 258208 57922 258278 57978
rect 258334 57922 258402 57978
rect 258458 57922 258528 57978
rect 258208 57888 258528 57922
rect 288928 58350 289248 58384
rect 288928 58294 288998 58350
rect 289054 58294 289122 58350
rect 289178 58294 289248 58350
rect 288928 58226 289248 58294
rect 288928 58170 288998 58226
rect 289054 58170 289122 58226
rect 289178 58170 289248 58226
rect 288928 58102 289248 58170
rect 288928 58046 288998 58102
rect 289054 58046 289122 58102
rect 289178 58046 289248 58102
rect 288928 57978 289248 58046
rect 288928 57922 288998 57978
rect 289054 57922 289122 57978
rect 289178 57922 289248 57978
rect 288928 57888 289248 57922
rect 319648 58350 319968 58384
rect 319648 58294 319718 58350
rect 319774 58294 319842 58350
rect 319898 58294 319968 58350
rect 319648 58226 319968 58294
rect 319648 58170 319718 58226
rect 319774 58170 319842 58226
rect 319898 58170 319968 58226
rect 319648 58102 319968 58170
rect 319648 58046 319718 58102
rect 319774 58046 319842 58102
rect 319898 58046 319968 58102
rect 319648 57978 319968 58046
rect 319648 57922 319718 57978
rect 319774 57922 319842 57978
rect 319898 57922 319968 57978
rect 319648 57888 319968 57922
rect 350368 58350 350688 58384
rect 350368 58294 350438 58350
rect 350494 58294 350562 58350
rect 350618 58294 350688 58350
rect 350368 58226 350688 58294
rect 350368 58170 350438 58226
rect 350494 58170 350562 58226
rect 350618 58170 350688 58226
rect 350368 58102 350688 58170
rect 350368 58046 350438 58102
rect 350494 58046 350562 58102
rect 350618 58046 350688 58102
rect 350368 57978 350688 58046
rect 350368 57922 350438 57978
rect 350494 57922 350562 57978
rect 350618 57922 350688 57978
rect 350368 57888 350688 57922
rect 381088 58350 381408 58384
rect 381088 58294 381158 58350
rect 381214 58294 381282 58350
rect 381338 58294 381408 58350
rect 381088 58226 381408 58294
rect 381088 58170 381158 58226
rect 381214 58170 381282 58226
rect 381338 58170 381408 58226
rect 381088 58102 381408 58170
rect 381088 58046 381158 58102
rect 381214 58046 381282 58102
rect 381338 58046 381408 58102
rect 381088 57978 381408 58046
rect 381088 57922 381158 57978
rect 381214 57922 381282 57978
rect 381338 57922 381408 57978
rect 381088 57888 381408 57922
rect 411808 58350 412128 58384
rect 411808 58294 411878 58350
rect 411934 58294 412002 58350
rect 412058 58294 412128 58350
rect 411808 58226 412128 58294
rect 411808 58170 411878 58226
rect 411934 58170 412002 58226
rect 412058 58170 412128 58226
rect 411808 58102 412128 58170
rect 411808 58046 411878 58102
rect 411934 58046 412002 58102
rect 412058 58046 412128 58102
rect 411808 57978 412128 58046
rect 411808 57922 411878 57978
rect 411934 57922 412002 57978
rect 412058 57922 412128 57978
rect 411808 57888 412128 57922
rect 442528 58350 442848 58384
rect 442528 58294 442598 58350
rect 442654 58294 442722 58350
rect 442778 58294 442848 58350
rect 442528 58226 442848 58294
rect 442528 58170 442598 58226
rect 442654 58170 442722 58226
rect 442778 58170 442848 58226
rect 442528 58102 442848 58170
rect 442528 58046 442598 58102
rect 442654 58046 442722 58102
rect 442778 58046 442848 58102
rect 442528 57978 442848 58046
rect 442528 57922 442598 57978
rect 442654 57922 442722 57978
rect 442778 57922 442848 57978
rect 442528 57888 442848 57922
rect 473248 58350 473568 58384
rect 473248 58294 473318 58350
rect 473374 58294 473442 58350
rect 473498 58294 473568 58350
rect 473248 58226 473568 58294
rect 473248 58170 473318 58226
rect 473374 58170 473442 58226
rect 473498 58170 473568 58226
rect 473248 58102 473568 58170
rect 473248 58046 473318 58102
rect 473374 58046 473442 58102
rect 473498 58046 473568 58102
rect 473248 57978 473568 58046
rect 473248 57922 473318 57978
rect 473374 57922 473442 57978
rect 473498 57922 473568 57978
rect 473248 57888 473568 57922
rect 503968 58350 504288 58384
rect 503968 58294 504038 58350
rect 504094 58294 504162 58350
rect 504218 58294 504288 58350
rect 503968 58226 504288 58294
rect 503968 58170 504038 58226
rect 504094 58170 504162 58226
rect 504218 58170 504288 58226
rect 503968 58102 504288 58170
rect 503968 58046 504038 58102
rect 504094 58046 504162 58102
rect 504218 58046 504288 58102
rect 503968 57978 504288 58046
rect 503968 57922 504038 57978
rect 504094 57922 504162 57978
rect 504218 57922 504288 57978
rect 503968 57888 504288 57922
rect 534688 58350 535008 58384
rect 534688 58294 534758 58350
rect 534814 58294 534882 58350
rect 534938 58294 535008 58350
rect 534688 58226 535008 58294
rect 534688 58170 534758 58226
rect 534814 58170 534882 58226
rect 534938 58170 535008 58226
rect 534688 58102 535008 58170
rect 534688 58046 534758 58102
rect 534814 58046 534882 58102
rect 534938 58046 535008 58102
rect 534688 57978 535008 58046
rect 534688 57922 534758 57978
rect 534814 57922 534882 57978
rect 534938 57922 535008 57978
rect 534688 57888 535008 57922
rect 565408 58350 565728 58384
rect 565408 58294 565478 58350
rect 565534 58294 565602 58350
rect 565658 58294 565728 58350
rect 565408 58226 565728 58294
rect 565408 58170 565478 58226
rect 565534 58170 565602 58226
rect 565658 58170 565728 58226
rect 565408 58102 565728 58170
rect 565408 58046 565478 58102
rect 565534 58046 565602 58102
rect 565658 58046 565728 58102
rect 565408 57978 565728 58046
rect 565408 57922 565478 57978
rect 565534 57922 565602 57978
rect 565658 57922 565728 57978
rect 565408 57888 565728 57922
rect 589098 58350 589718 75922
rect 589098 58294 589194 58350
rect 589250 58294 589318 58350
rect 589374 58294 589442 58350
rect 589498 58294 589566 58350
rect 589622 58294 589718 58350
rect 589098 58226 589718 58294
rect 589098 58170 589194 58226
rect 589250 58170 589318 58226
rect 589374 58170 589442 58226
rect 589498 58170 589566 58226
rect 589622 58170 589718 58226
rect 589098 58102 589718 58170
rect 589098 58046 589194 58102
rect 589250 58046 589318 58102
rect 589374 58046 589442 58102
rect 589498 58046 589566 58102
rect 589622 58046 589718 58102
rect 589098 57978 589718 58046
rect 589098 57922 589194 57978
rect 589250 57922 589318 57978
rect 589374 57922 589442 57978
rect 589498 57922 589566 57978
rect 589622 57922 589718 57978
rect 27808 46350 28128 46384
rect 27808 46294 27878 46350
rect 27934 46294 28002 46350
rect 28058 46294 28128 46350
rect 27808 46226 28128 46294
rect 27808 46170 27878 46226
rect 27934 46170 28002 46226
rect 28058 46170 28128 46226
rect 27808 46102 28128 46170
rect 27808 46046 27878 46102
rect 27934 46046 28002 46102
rect 28058 46046 28128 46102
rect 27808 45978 28128 46046
rect 27808 45922 27878 45978
rect 27934 45922 28002 45978
rect 28058 45922 28128 45978
rect 27808 45888 28128 45922
rect 58528 46350 58848 46384
rect 58528 46294 58598 46350
rect 58654 46294 58722 46350
rect 58778 46294 58848 46350
rect 58528 46226 58848 46294
rect 58528 46170 58598 46226
rect 58654 46170 58722 46226
rect 58778 46170 58848 46226
rect 58528 46102 58848 46170
rect 58528 46046 58598 46102
rect 58654 46046 58722 46102
rect 58778 46046 58848 46102
rect 58528 45978 58848 46046
rect 58528 45922 58598 45978
rect 58654 45922 58722 45978
rect 58778 45922 58848 45978
rect 58528 45888 58848 45922
rect 89248 46350 89568 46384
rect 89248 46294 89318 46350
rect 89374 46294 89442 46350
rect 89498 46294 89568 46350
rect 89248 46226 89568 46294
rect 89248 46170 89318 46226
rect 89374 46170 89442 46226
rect 89498 46170 89568 46226
rect 89248 46102 89568 46170
rect 89248 46046 89318 46102
rect 89374 46046 89442 46102
rect 89498 46046 89568 46102
rect 89248 45978 89568 46046
rect 89248 45922 89318 45978
rect 89374 45922 89442 45978
rect 89498 45922 89568 45978
rect 89248 45888 89568 45922
rect 119968 46350 120288 46384
rect 119968 46294 120038 46350
rect 120094 46294 120162 46350
rect 120218 46294 120288 46350
rect 119968 46226 120288 46294
rect 119968 46170 120038 46226
rect 120094 46170 120162 46226
rect 120218 46170 120288 46226
rect 119968 46102 120288 46170
rect 119968 46046 120038 46102
rect 120094 46046 120162 46102
rect 120218 46046 120288 46102
rect 119968 45978 120288 46046
rect 119968 45922 120038 45978
rect 120094 45922 120162 45978
rect 120218 45922 120288 45978
rect 119968 45888 120288 45922
rect 150688 46350 151008 46384
rect 150688 46294 150758 46350
rect 150814 46294 150882 46350
rect 150938 46294 151008 46350
rect 150688 46226 151008 46294
rect 150688 46170 150758 46226
rect 150814 46170 150882 46226
rect 150938 46170 151008 46226
rect 150688 46102 151008 46170
rect 150688 46046 150758 46102
rect 150814 46046 150882 46102
rect 150938 46046 151008 46102
rect 150688 45978 151008 46046
rect 150688 45922 150758 45978
rect 150814 45922 150882 45978
rect 150938 45922 151008 45978
rect 150688 45888 151008 45922
rect 181408 46350 181728 46384
rect 181408 46294 181478 46350
rect 181534 46294 181602 46350
rect 181658 46294 181728 46350
rect 181408 46226 181728 46294
rect 181408 46170 181478 46226
rect 181534 46170 181602 46226
rect 181658 46170 181728 46226
rect 181408 46102 181728 46170
rect 181408 46046 181478 46102
rect 181534 46046 181602 46102
rect 181658 46046 181728 46102
rect 181408 45978 181728 46046
rect 181408 45922 181478 45978
rect 181534 45922 181602 45978
rect 181658 45922 181728 45978
rect 181408 45888 181728 45922
rect 212128 46350 212448 46384
rect 212128 46294 212198 46350
rect 212254 46294 212322 46350
rect 212378 46294 212448 46350
rect 212128 46226 212448 46294
rect 212128 46170 212198 46226
rect 212254 46170 212322 46226
rect 212378 46170 212448 46226
rect 212128 46102 212448 46170
rect 212128 46046 212198 46102
rect 212254 46046 212322 46102
rect 212378 46046 212448 46102
rect 212128 45978 212448 46046
rect 212128 45922 212198 45978
rect 212254 45922 212322 45978
rect 212378 45922 212448 45978
rect 212128 45888 212448 45922
rect 242848 46350 243168 46384
rect 242848 46294 242918 46350
rect 242974 46294 243042 46350
rect 243098 46294 243168 46350
rect 242848 46226 243168 46294
rect 242848 46170 242918 46226
rect 242974 46170 243042 46226
rect 243098 46170 243168 46226
rect 242848 46102 243168 46170
rect 242848 46046 242918 46102
rect 242974 46046 243042 46102
rect 243098 46046 243168 46102
rect 242848 45978 243168 46046
rect 242848 45922 242918 45978
rect 242974 45922 243042 45978
rect 243098 45922 243168 45978
rect 242848 45888 243168 45922
rect 273568 46350 273888 46384
rect 273568 46294 273638 46350
rect 273694 46294 273762 46350
rect 273818 46294 273888 46350
rect 273568 46226 273888 46294
rect 273568 46170 273638 46226
rect 273694 46170 273762 46226
rect 273818 46170 273888 46226
rect 273568 46102 273888 46170
rect 273568 46046 273638 46102
rect 273694 46046 273762 46102
rect 273818 46046 273888 46102
rect 273568 45978 273888 46046
rect 273568 45922 273638 45978
rect 273694 45922 273762 45978
rect 273818 45922 273888 45978
rect 273568 45888 273888 45922
rect 304288 46350 304608 46384
rect 304288 46294 304358 46350
rect 304414 46294 304482 46350
rect 304538 46294 304608 46350
rect 304288 46226 304608 46294
rect 304288 46170 304358 46226
rect 304414 46170 304482 46226
rect 304538 46170 304608 46226
rect 304288 46102 304608 46170
rect 304288 46046 304358 46102
rect 304414 46046 304482 46102
rect 304538 46046 304608 46102
rect 304288 45978 304608 46046
rect 304288 45922 304358 45978
rect 304414 45922 304482 45978
rect 304538 45922 304608 45978
rect 304288 45888 304608 45922
rect 335008 46350 335328 46384
rect 335008 46294 335078 46350
rect 335134 46294 335202 46350
rect 335258 46294 335328 46350
rect 335008 46226 335328 46294
rect 335008 46170 335078 46226
rect 335134 46170 335202 46226
rect 335258 46170 335328 46226
rect 335008 46102 335328 46170
rect 335008 46046 335078 46102
rect 335134 46046 335202 46102
rect 335258 46046 335328 46102
rect 335008 45978 335328 46046
rect 335008 45922 335078 45978
rect 335134 45922 335202 45978
rect 335258 45922 335328 45978
rect 335008 45888 335328 45922
rect 365728 46350 366048 46384
rect 365728 46294 365798 46350
rect 365854 46294 365922 46350
rect 365978 46294 366048 46350
rect 365728 46226 366048 46294
rect 365728 46170 365798 46226
rect 365854 46170 365922 46226
rect 365978 46170 366048 46226
rect 365728 46102 366048 46170
rect 365728 46046 365798 46102
rect 365854 46046 365922 46102
rect 365978 46046 366048 46102
rect 365728 45978 366048 46046
rect 365728 45922 365798 45978
rect 365854 45922 365922 45978
rect 365978 45922 366048 45978
rect 365728 45888 366048 45922
rect 396448 46350 396768 46384
rect 396448 46294 396518 46350
rect 396574 46294 396642 46350
rect 396698 46294 396768 46350
rect 396448 46226 396768 46294
rect 396448 46170 396518 46226
rect 396574 46170 396642 46226
rect 396698 46170 396768 46226
rect 396448 46102 396768 46170
rect 396448 46046 396518 46102
rect 396574 46046 396642 46102
rect 396698 46046 396768 46102
rect 396448 45978 396768 46046
rect 396448 45922 396518 45978
rect 396574 45922 396642 45978
rect 396698 45922 396768 45978
rect 396448 45888 396768 45922
rect 427168 46350 427488 46384
rect 427168 46294 427238 46350
rect 427294 46294 427362 46350
rect 427418 46294 427488 46350
rect 427168 46226 427488 46294
rect 427168 46170 427238 46226
rect 427294 46170 427362 46226
rect 427418 46170 427488 46226
rect 427168 46102 427488 46170
rect 427168 46046 427238 46102
rect 427294 46046 427362 46102
rect 427418 46046 427488 46102
rect 427168 45978 427488 46046
rect 427168 45922 427238 45978
rect 427294 45922 427362 45978
rect 427418 45922 427488 45978
rect 427168 45888 427488 45922
rect 457888 46350 458208 46384
rect 457888 46294 457958 46350
rect 458014 46294 458082 46350
rect 458138 46294 458208 46350
rect 457888 46226 458208 46294
rect 457888 46170 457958 46226
rect 458014 46170 458082 46226
rect 458138 46170 458208 46226
rect 457888 46102 458208 46170
rect 457888 46046 457958 46102
rect 458014 46046 458082 46102
rect 458138 46046 458208 46102
rect 457888 45978 458208 46046
rect 457888 45922 457958 45978
rect 458014 45922 458082 45978
rect 458138 45922 458208 45978
rect 457888 45888 458208 45922
rect 488608 46350 488928 46384
rect 488608 46294 488678 46350
rect 488734 46294 488802 46350
rect 488858 46294 488928 46350
rect 488608 46226 488928 46294
rect 488608 46170 488678 46226
rect 488734 46170 488802 46226
rect 488858 46170 488928 46226
rect 488608 46102 488928 46170
rect 488608 46046 488678 46102
rect 488734 46046 488802 46102
rect 488858 46046 488928 46102
rect 488608 45978 488928 46046
rect 488608 45922 488678 45978
rect 488734 45922 488802 45978
rect 488858 45922 488928 45978
rect 488608 45888 488928 45922
rect 519328 46350 519648 46384
rect 519328 46294 519398 46350
rect 519454 46294 519522 46350
rect 519578 46294 519648 46350
rect 519328 46226 519648 46294
rect 519328 46170 519398 46226
rect 519454 46170 519522 46226
rect 519578 46170 519648 46226
rect 519328 46102 519648 46170
rect 519328 46046 519398 46102
rect 519454 46046 519522 46102
rect 519578 46046 519648 46102
rect 519328 45978 519648 46046
rect 519328 45922 519398 45978
rect 519454 45922 519522 45978
rect 519578 45922 519648 45978
rect 519328 45888 519648 45922
rect 550048 46350 550368 46384
rect 550048 46294 550118 46350
rect 550174 46294 550242 46350
rect 550298 46294 550368 46350
rect 550048 46226 550368 46294
rect 550048 46170 550118 46226
rect 550174 46170 550242 46226
rect 550298 46170 550368 46226
rect 550048 46102 550368 46170
rect 550048 46046 550118 46102
rect 550174 46046 550242 46102
rect 550298 46046 550368 46102
rect 550048 45978 550368 46046
rect 550048 45922 550118 45978
rect 550174 45922 550242 45978
rect 550298 45922 550368 45978
rect 550048 45888 550368 45922
rect 5418 40294 5514 40350
rect 5570 40294 5638 40350
rect 5694 40294 5762 40350
rect 5818 40294 5886 40350
rect 5942 40294 6038 40350
rect 5418 40226 6038 40294
rect 5418 40170 5514 40226
rect 5570 40170 5638 40226
rect 5694 40170 5762 40226
rect 5818 40170 5886 40226
rect 5942 40170 6038 40226
rect 5418 40102 6038 40170
rect 5418 40046 5514 40102
rect 5570 40046 5638 40102
rect 5694 40046 5762 40102
rect 5818 40046 5886 40102
rect 5942 40046 6038 40102
rect 5418 39978 6038 40046
rect 5418 39922 5514 39978
rect 5570 39922 5638 39978
rect 5694 39922 5762 39978
rect 5818 39922 5886 39978
rect 5942 39922 6038 39978
rect 4060 38724 4116 38734
rect 4060 36932 4116 38668
rect 4060 36866 4116 36876
rect 4172 28196 4228 28206
rect 4172 22932 4228 28140
rect 4172 22866 4228 22876
rect -956 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 -336 22350
rect -956 22226 -336 22294
rect -956 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 -336 22226
rect -956 22102 -336 22170
rect -956 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 -336 22102
rect -956 21978 -336 22046
rect -956 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 -336 21978
rect -956 4350 -336 21922
rect -956 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 -336 4350
rect -956 4226 -336 4294
rect -956 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 -336 4226
rect -956 4102 -336 4170
rect -956 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 -336 4102
rect -956 3978 -336 4046
rect -956 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 -336 3978
rect -956 -160 -336 3922
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 -336 -160
rect -956 -284 -336 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 -336 -284
rect -956 -408 -336 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 -336 -408
rect -956 -532 -336 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 -336 -532
rect -956 -684 -336 -588
rect 5418 22350 6038 39922
rect 12448 40350 12768 40384
rect 12448 40294 12518 40350
rect 12574 40294 12642 40350
rect 12698 40294 12768 40350
rect 12448 40226 12768 40294
rect 12448 40170 12518 40226
rect 12574 40170 12642 40226
rect 12698 40170 12768 40226
rect 12448 40102 12768 40170
rect 12448 40046 12518 40102
rect 12574 40046 12642 40102
rect 12698 40046 12768 40102
rect 12448 39978 12768 40046
rect 12448 39922 12518 39978
rect 12574 39922 12642 39978
rect 12698 39922 12768 39978
rect 12448 39888 12768 39922
rect 43168 40350 43488 40384
rect 43168 40294 43238 40350
rect 43294 40294 43362 40350
rect 43418 40294 43488 40350
rect 43168 40226 43488 40294
rect 43168 40170 43238 40226
rect 43294 40170 43362 40226
rect 43418 40170 43488 40226
rect 43168 40102 43488 40170
rect 43168 40046 43238 40102
rect 43294 40046 43362 40102
rect 43418 40046 43488 40102
rect 43168 39978 43488 40046
rect 43168 39922 43238 39978
rect 43294 39922 43362 39978
rect 43418 39922 43488 39978
rect 43168 39888 43488 39922
rect 73888 40350 74208 40384
rect 73888 40294 73958 40350
rect 74014 40294 74082 40350
rect 74138 40294 74208 40350
rect 73888 40226 74208 40294
rect 73888 40170 73958 40226
rect 74014 40170 74082 40226
rect 74138 40170 74208 40226
rect 73888 40102 74208 40170
rect 73888 40046 73958 40102
rect 74014 40046 74082 40102
rect 74138 40046 74208 40102
rect 73888 39978 74208 40046
rect 73888 39922 73958 39978
rect 74014 39922 74082 39978
rect 74138 39922 74208 39978
rect 73888 39888 74208 39922
rect 104608 40350 104928 40384
rect 104608 40294 104678 40350
rect 104734 40294 104802 40350
rect 104858 40294 104928 40350
rect 104608 40226 104928 40294
rect 104608 40170 104678 40226
rect 104734 40170 104802 40226
rect 104858 40170 104928 40226
rect 104608 40102 104928 40170
rect 104608 40046 104678 40102
rect 104734 40046 104802 40102
rect 104858 40046 104928 40102
rect 104608 39978 104928 40046
rect 104608 39922 104678 39978
rect 104734 39922 104802 39978
rect 104858 39922 104928 39978
rect 104608 39888 104928 39922
rect 135328 40350 135648 40384
rect 135328 40294 135398 40350
rect 135454 40294 135522 40350
rect 135578 40294 135648 40350
rect 135328 40226 135648 40294
rect 135328 40170 135398 40226
rect 135454 40170 135522 40226
rect 135578 40170 135648 40226
rect 135328 40102 135648 40170
rect 135328 40046 135398 40102
rect 135454 40046 135522 40102
rect 135578 40046 135648 40102
rect 135328 39978 135648 40046
rect 135328 39922 135398 39978
rect 135454 39922 135522 39978
rect 135578 39922 135648 39978
rect 135328 39888 135648 39922
rect 166048 40350 166368 40384
rect 166048 40294 166118 40350
rect 166174 40294 166242 40350
rect 166298 40294 166368 40350
rect 166048 40226 166368 40294
rect 166048 40170 166118 40226
rect 166174 40170 166242 40226
rect 166298 40170 166368 40226
rect 166048 40102 166368 40170
rect 166048 40046 166118 40102
rect 166174 40046 166242 40102
rect 166298 40046 166368 40102
rect 166048 39978 166368 40046
rect 166048 39922 166118 39978
rect 166174 39922 166242 39978
rect 166298 39922 166368 39978
rect 166048 39888 166368 39922
rect 196768 40350 197088 40384
rect 196768 40294 196838 40350
rect 196894 40294 196962 40350
rect 197018 40294 197088 40350
rect 196768 40226 197088 40294
rect 196768 40170 196838 40226
rect 196894 40170 196962 40226
rect 197018 40170 197088 40226
rect 196768 40102 197088 40170
rect 196768 40046 196838 40102
rect 196894 40046 196962 40102
rect 197018 40046 197088 40102
rect 196768 39978 197088 40046
rect 196768 39922 196838 39978
rect 196894 39922 196962 39978
rect 197018 39922 197088 39978
rect 196768 39888 197088 39922
rect 227488 40350 227808 40384
rect 227488 40294 227558 40350
rect 227614 40294 227682 40350
rect 227738 40294 227808 40350
rect 227488 40226 227808 40294
rect 227488 40170 227558 40226
rect 227614 40170 227682 40226
rect 227738 40170 227808 40226
rect 227488 40102 227808 40170
rect 227488 40046 227558 40102
rect 227614 40046 227682 40102
rect 227738 40046 227808 40102
rect 227488 39978 227808 40046
rect 227488 39922 227558 39978
rect 227614 39922 227682 39978
rect 227738 39922 227808 39978
rect 227488 39888 227808 39922
rect 258208 40350 258528 40384
rect 258208 40294 258278 40350
rect 258334 40294 258402 40350
rect 258458 40294 258528 40350
rect 258208 40226 258528 40294
rect 258208 40170 258278 40226
rect 258334 40170 258402 40226
rect 258458 40170 258528 40226
rect 258208 40102 258528 40170
rect 258208 40046 258278 40102
rect 258334 40046 258402 40102
rect 258458 40046 258528 40102
rect 258208 39978 258528 40046
rect 258208 39922 258278 39978
rect 258334 39922 258402 39978
rect 258458 39922 258528 39978
rect 258208 39888 258528 39922
rect 288928 40350 289248 40384
rect 288928 40294 288998 40350
rect 289054 40294 289122 40350
rect 289178 40294 289248 40350
rect 288928 40226 289248 40294
rect 288928 40170 288998 40226
rect 289054 40170 289122 40226
rect 289178 40170 289248 40226
rect 288928 40102 289248 40170
rect 288928 40046 288998 40102
rect 289054 40046 289122 40102
rect 289178 40046 289248 40102
rect 288928 39978 289248 40046
rect 288928 39922 288998 39978
rect 289054 39922 289122 39978
rect 289178 39922 289248 39978
rect 288928 39888 289248 39922
rect 319648 40350 319968 40384
rect 319648 40294 319718 40350
rect 319774 40294 319842 40350
rect 319898 40294 319968 40350
rect 319648 40226 319968 40294
rect 319648 40170 319718 40226
rect 319774 40170 319842 40226
rect 319898 40170 319968 40226
rect 319648 40102 319968 40170
rect 319648 40046 319718 40102
rect 319774 40046 319842 40102
rect 319898 40046 319968 40102
rect 319648 39978 319968 40046
rect 319648 39922 319718 39978
rect 319774 39922 319842 39978
rect 319898 39922 319968 39978
rect 319648 39888 319968 39922
rect 350368 40350 350688 40384
rect 350368 40294 350438 40350
rect 350494 40294 350562 40350
rect 350618 40294 350688 40350
rect 350368 40226 350688 40294
rect 350368 40170 350438 40226
rect 350494 40170 350562 40226
rect 350618 40170 350688 40226
rect 350368 40102 350688 40170
rect 350368 40046 350438 40102
rect 350494 40046 350562 40102
rect 350618 40046 350688 40102
rect 350368 39978 350688 40046
rect 350368 39922 350438 39978
rect 350494 39922 350562 39978
rect 350618 39922 350688 39978
rect 350368 39888 350688 39922
rect 381088 40350 381408 40384
rect 381088 40294 381158 40350
rect 381214 40294 381282 40350
rect 381338 40294 381408 40350
rect 381088 40226 381408 40294
rect 381088 40170 381158 40226
rect 381214 40170 381282 40226
rect 381338 40170 381408 40226
rect 381088 40102 381408 40170
rect 381088 40046 381158 40102
rect 381214 40046 381282 40102
rect 381338 40046 381408 40102
rect 381088 39978 381408 40046
rect 381088 39922 381158 39978
rect 381214 39922 381282 39978
rect 381338 39922 381408 39978
rect 381088 39888 381408 39922
rect 411808 40350 412128 40384
rect 411808 40294 411878 40350
rect 411934 40294 412002 40350
rect 412058 40294 412128 40350
rect 411808 40226 412128 40294
rect 411808 40170 411878 40226
rect 411934 40170 412002 40226
rect 412058 40170 412128 40226
rect 411808 40102 412128 40170
rect 411808 40046 411878 40102
rect 411934 40046 412002 40102
rect 412058 40046 412128 40102
rect 411808 39978 412128 40046
rect 411808 39922 411878 39978
rect 411934 39922 412002 39978
rect 412058 39922 412128 39978
rect 411808 39888 412128 39922
rect 442528 40350 442848 40384
rect 442528 40294 442598 40350
rect 442654 40294 442722 40350
rect 442778 40294 442848 40350
rect 442528 40226 442848 40294
rect 442528 40170 442598 40226
rect 442654 40170 442722 40226
rect 442778 40170 442848 40226
rect 442528 40102 442848 40170
rect 442528 40046 442598 40102
rect 442654 40046 442722 40102
rect 442778 40046 442848 40102
rect 442528 39978 442848 40046
rect 442528 39922 442598 39978
rect 442654 39922 442722 39978
rect 442778 39922 442848 39978
rect 442528 39888 442848 39922
rect 473248 40350 473568 40384
rect 473248 40294 473318 40350
rect 473374 40294 473442 40350
rect 473498 40294 473568 40350
rect 473248 40226 473568 40294
rect 473248 40170 473318 40226
rect 473374 40170 473442 40226
rect 473498 40170 473568 40226
rect 473248 40102 473568 40170
rect 473248 40046 473318 40102
rect 473374 40046 473442 40102
rect 473498 40046 473568 40102
rect 473248 39978 473568 40046
rect 473248 39922 473318 39978
rect 473374 39922 473442 39978
rect 473498 39922 473568 39978
rect 473248 39888 473568 39922
rect 503968 40350 504288 40384
rect 503968 40294 504038 40350
rect 504094 40294 504162 40350
rect 504218 40294 504288 40350
rect 503968 40226 504288 40294
rect 503968 40170 504038 40226
rect 504094 40170 504162 40226
rect 504218 40170 504288 40226
rect 503968 40102 504288 40170
rect 503968 40046 504038 40102
rect 504094 40046 504162 40102
rect 504218 40046 504288 40102
rect 503968 39978 504288 40046
rect 503968 39922 504038 39978
rect 504094 39922 504162 39978
rect 504218 39922 504288 39978
rect 503968 39888 504288 39922
rect 534688 40350 535008 40384
rect 534688 40294 534758 40350
rect 534814 40294 534882 40350
rect 534938 40294 535008 40350
rect 534688 40226 535008 40294
rect 534688 40170 534758 40226
rect 534814 40170 534882 40226
rect 534938 40170 535008 40226
rect 534688 40102 535008 40170
rect 534688 40046 534758 40102
rect 534814 40046 534882 40102
rect 534938 40046 535008 40102
rect 534688 39978 535008 40046
rect 534688 39922 534758 39978
rect 534814 39922 534882 39978
rect 534938 39922 535008 39978
rect 534688 39888 535008 39922
rect 565408 40350 565728 40384
rect 565408 40294 565478 40350
rect 565534 40294 565602 40350
rect 565658 40294 565728 40350
rect 565408 40226 565728 40294
rect 565408 40170 565478 40226
rect 565534 40170 565602 40226
rect 565658 40170 565728 40226
rect 565408 40102 565728 40170
rect 565408 40046 565478 40102
rect 565534 40046 565602 40102
rect 565658 40046 565728 40102
rect 565408 39978 565728 40046
rect 565408 39922 565478 39978
rect 565534 39922 565602 39978
rect 565658 39922 565728 39978
rect 565408 39888 565728 39922
rect 589098 40350 589718 57922
rect 592818 64350 593438 81922
rect 592818 64294 592914 64350
rect 592970 64294 593038 64350
rect 593094 64294 593162 64350
rect 593218 64294 593286 64350
rect 593342 64294 593438 64350
rect 592818 64226 593438 64294
rect 592818 64170 592914 64226
rect 592970 64170 593038 64226
rect 593094 64170 593162 64226
rect 593218 64170 593286 64226
rect 593342 64170 593438 64226
rect 592818 64102 593438 64170
rect 592818 64046 592914 64102
rect 592970 64046 593038 64102
rect 593094 64046 593162 64102
rect 593218 64046 593286 64102
rect 593342 64046 593438 64102
rect 592818 63978 593438 64046
rect 592818 63922 592914 63978
rect 592970 63922 593038 63978
rect 593094 63922 593162 63978
rect 593218 63922 593286 63978
rect 593342 63922 593438 63978
rect 590492 49476 590548 49486
rect 590492 47012 590548 49420
rect 590492 46946 590548 46956
rect 589098 40294 589194 40350
rect 589250 40294 589318 40350
rect 589374 40294 589442 40350
rect 589498 40294 589566 40350
rect 589622 40294 589718 40350
rect 589098 40226 589718 40294
rect 589098 40170 589194 40226
rect 589250 40170 589318 40226
rect 589374 40170 589442 40226
rect 589498 40170 589566 40226
rect 589622 40170 589718 40226
rect 589098 40102 589718 40170
rect 589098 40046 589194 40102
rect 589250 40046 589318 40102
rect 589374 40046 589442 40102
rect 589498 40046 589566 40102
rect 589622 40046 589718 40102
rect 589098 39978 589718 40046
rect 589098 39922 589194 39978
rect 589250 39922 589318 39978
rect 589374 39922 589442 39978
rect 589498 39922 589566 39978
rect 589622 39922 589718 39978
rect 588812 38724 588868 38734
rect 588812 33796 588868 38668
rect 588812 33730 588868 33740
rect 27808 28350 28128 28384
rect 27808 28294 27878 28350
rect 27934 28294 28002 28350
rect 28058 28294 28128 28350
rect 27808 28226 28128 28294
rect 27808 28170 27878 28226
rect 27934 28170 28002 28226
rect 28058 28170 28128 28226
rect 27808 28102 28128 28170
rect 27808 28046 27878 28102
rect 27934 28046 28002 28102
rect 28058 28046 28128 28102
rect 27808 27978 28128 28046
rect 27808 27922 27878 27978
rect 27934 27922 28002 27978
rect 28058 27922 28128 27978
rect 27808 27888 28128 27922
rect 58528 28350 58848 28384
rect 58528 28294 58598 28350
rect 58654 28294 58722 28350
rect 58778 28294 58848 28350
rect 58528 28226 58848 28294
rect 58528 28170 58598 28226
rect 58654 28170 58722 28226
rect 58778 28170 58848 28226
rect 58528 28102 58848 28170
rect 58528 28046 58598 28102
rect 58654 28046 58722 28102
rect 58778 28046 58848 28102
rect 58528 27978 58848 28046
rect 58528 27922 58598 27978
rect 58654 27922 58722 27978
rect 58778 27922 58848 27978
rect 58528 27888 58848 27922
rect 89248 28350 89568 28384
rect 89248 28294 89318 28350
rect 89374 28294 89442 28350
rect 89498 28294 89568 28350
rect 89248 28226 89568 28294
rect 89248 28170 89318 28226
rect 89374 28170 89442 28226
rect 89498 28170 89568 28226
rect 89248 28102 89568 28170
rect 89248 28046 89318 28102
rect 89374 28046 89442 28102
rect 89498 28046 89568 28102
rect 89248 27978 89568 28046
rect 89248 27922 89318 27978
rect 89374 27922 89442 27978
rect 89498 27922 89568 27978
rect 89248 27888 89568 27922
rect 119968 28350 120288 28384
rect 119968 28294 120038 28350
rect 120094 28294 120162 28350
rect 120218 28294 120288 28350
rect 119968 28226 120288 28294
rect 119968 28170 120038 28226
rect 120094 28170 120162 28226
rect 120218 28170 120288 28226
rect 119968 28102 120288 28170
rect 119968 28046 120038 28102
rect 120094 28046 120162 28102
rect 120218 28046 120288 28102
rect 119968 27978 120288 28046
rect 119968 27922 120038 27978
rect 120094 27922 120162 27978
rect 120218 27922 120288 27978
rect 119968 27888 120288 27922
rect 150688 28350 151008 28384
rect 150688 28294 150758 28350
rect 150814 28294 150882 28350
rect 150938 28294 151008 28350
rect 150688 28226 151008 28294
rect 150688 28170 150758 28226
rect 150814 28170 150882 28226
rect 150938 28170 151008 28226
rect 150688 28102 151008 28170
rect 150688 28046 150758 28102
rect 150814 28046 150882 28102
rect 150938 28046 151008 28102
rect 150688 27978 151008 28046
rect 150688 27922 150758 27978
rect 150814 27922 150882 27978
rect 150938 27922 151008 27978
rect 150688 27888 151008 27922
rect 181408 28350 181728 28384
rect 181408 28294 181478 28350
rect 181534 28294 181602 28350
rect 181658 28294 181728 28350
rect 181408 28226 181728 28294
rect 181408 28170 181478 28226
rect 181534 28170 181602 28226
rect 181658 28170 181728 28226
rect 181408 28102 181728 28170
rect 181408 28046 181478 28102
rect 181534 28046 181602 28102
rect 181658 28046 181728 28102
rect 181408 27978 181728 28046
rect 181408 27922 181478 27978
rect 181534 27922 181602 27978
rect 181658 27922 181728 27978
rect 181408 27888 181728 27922
rect 212128 28350 212448 28384
rect 212128 28294 212198 28350
rect 212254 28294 212322 28350
rect 212378 28294 212448 28350
rect 212128 28226 212448 28294
rect 212128 28170 212198 28226
rect 212254 28170 212322 28226
rect 212378 28170 212448 28226
rect 212128 28102 212448 28170
rect 212128 28046 212198 28102
rect 212254 28046 212322 28102
rect 212378 28046 212448 28102
rect 212128 27978 212448 28046
rect 212128 27922 212198 27978
rect 212254 27922 212322 27978
rect 212378 27922 212448 27978
rect 212128 27888 212448 27922
rect 242848 28350 243168 28384
rect 242848 28294 242918 28350
rect 242974 28294 243042 28350
rect 243098 28294 243168 28350
rect 242848 28226 243168 28294
rect 242848 28170 242918 28226
rect 242974 28170 243042 28226
rect 243098 28170 243168 28226
rect 242848 28102 243168 28170
rect 242848 28046 242918 28102
rect 242974 28046 243042 28102
rect 243098 28046 243168 28102
rect 242848 27978 243168 28046
rect 242848 27922 242918 27978
rect 242974 27922 243042 27978
rect 243098 27922 243168 27978
rect 242848 27888 243168 27922
rect 273568 28350 273888 28384
rect 273568 28294 273638 28350
rect 273694 28294 273762 28350
rect 273818 28294 273888 28350
rect 273568 28226 273888 28294
rect 273568 28170 273638 28226
rect 273694 28170 273762 28226
rect 273818 28170 273888 28226
rect 273568 28102 273888 28170
rect 273568 28046 273638 28102
rect 273694 28046 273762 28102
rect 273818 28046 273888 28102
rect 273568 27978 273888 28046
rect 273568 27922 273638 27978
rect 273694 27922 273762 27978
rect 273818 27922 273888 27978
rect 273568 27888 273888 27922
rect 304288 28350 304608 28384
rect 304288 28294 304358 28350
rect 304414 28294 304482 28350
rect 304538 28294 304608 28350
rect 304288 28226 304608 28294
rect 304288 28170 304358 28226
rect 304414 28170 304482 28226
rect 304538 28170 304608 28226
rect 304288 28102 304608 28170
rect 304288 28046 304358 28102
rect 304414 28046 304482 28102
rect 304538 28046 304608 28102
rect 304288 27978 304608 28046
rect 304288 27922 304358 27978
rect 304414 27922 304482 27978
rect 304538 27922 304608 27978
rect 304288 27888 304608 27922
rect 335008 28350 335328 28384
rect 335008 28294 335078 28350
rect 335134 28294 335202 28350
rect 335258 28294 335328 28350
rect 335008 28226 335328 28294
rect 335008 28170 335078 28226
rect 335134 28170 335202 28226
rect 335258 28170 335328 28226
rect 335008 28102 335328 28170
rect 335008 28046 335078 28102
rect 335134 28046 335202 28102
rect 335258 28046 335328 28102
rect 335008 27978 335328 28046
rect 335008 27922 335078 27978
rect 335134 27922 335202 27978
rect 335258 27922 335328 27978
rect 335008 27888 335328 27922
rect 365728 28350 366048 28384
rect 365728 28294 365798 28350
rect 365854 28294 365922 28350
rect 365978 28294 366048 28350
rect 365728 28226 366048 28294
rect 365728 28170 365798 28226
rect 365854 28170 365922 28226
rect 365978 28170 366048 28226
rect 365728 28102 366048 28170
rect 365728 28046 365798 28102
rect 365854 28046 365922 28102
rect 365978 28046 366048 28102
rect 365728 27978 366048 28046
rect 365728 27922 365798 27978
rect 365854 27922 365922 27978
rect 365978 27922 366048 27978
rect 365728 27888 366048 27922
rect 396448 28350 396768 28384
rect 396448 28294 396518 28350
rect 396574 28294 396642 28350
rect 396698 28294 396768 28350
rect 396448 28226 396768 28294
rect 396448 28170 396518 28226
rect 396574 28170 396642 28226
rect 396698 28170 396768 28226
rect 396448 28102 396768 28170
rect 396448 28046 396518 28102
rect 396574 28046 396642 28102
rect 396698 28046 396768 28102
rect 396448 27978 396768 28046
rect 396448 27922 396518 27978
rect 396574 27922 396642 27978
rect 396698 27922 396768 27978
rect 396448 27888 396768 27922
rect 427168 28350 427488 28384
rect 427168 28294 427238 28350
rect 427294 28294 427362 28350
rect 427418 28294 427488 28350
rect 427168 28226 427488 28294
rect 427168 28170 427238 28226
rect 427294 28170 427362 28226
rect 427418 28170 427488 28226
rect 427168 28102 427488 28170
rect 427168 28046 427238 28102
rect 427294 28046 427362 28102
rect 427418 28046 427488 28102
rect 427168 27978 427488 28046
rect 427168 27922 427238 27978
rect 427294 27922 427362 27978
rect 427418 27922 427488 27978
rect 427168 27888 427488 27922
rect 457888 28350 458208 28384
rect 457888 28294 457958 28350
rect 458014 28294 458082 28350
rect 458138 28294 458208 28350
rect 457888 28226 458208 28294
rect 457888 28170 457958 28226
rect 458014 28170 458082 28226
rect 458138 28170 458208 28226
rect 457888 28102 458208 28170
rect 457888 28046 457958 28102
rect 458014 28046 458082 28102
rect 458138 28046 458208 28102
rect 457888 27978 458208 28046
rect 457888 27922 457958 27978
rect 458014 27922 458082 27978
rect 458138 27922 458208 27978
rect 457888 27888 458208 27922
rect 488608 28350 488928 28384
rect 488608 28294 488678 28350
rect 488734 28294 488802 28350
rect 488858 28294 488928 28350
rect 488608 28226 488928 28294
rect 488608 28170 488678 28226
rect 488734 28170 488802 28226
rect 488858 28170 488928 28226
rect 488608 28102 488928 28170
rect 488608 28046 488678 28102
rect 488734 28046 488802 28102
rect 488858 28046 488928 28102
rect 488608 27978 488928 28046
rect 488608 27922 488678 27978
rect 488734 27922 488802 27978
rect 488858 27922 488928 27978
rect 488608 27888 488928 27922
rect 519328 28350 519648 28384
rect 519328 28294 519398 28350
rect 519454 28294 519522 28350
rect 519578 28294 519648 28350
rect 519328 28226 519648 28294
rect 519328 28170 519398 28226
rect 519454 28170 519522 28226
rect 519578 28170 519648 28226
rect 519328 28102 519648 28170
rect 519328 28046 519398 28102
rect 519454 28046 519522 28102
rect 519578 28046 519648 28102
rect 519328 27978 519648 28046
rect 519328 27922 519398 27978
rect 519454 27922 519522 27978
rect 519578 27922 519648 27978
rect 519328 27888 519648 27922
rect 550048 28350 550368 28384
rect 550048 28294 550118 28350
rect 550174 28294 550242 28350
rect 550298 28294 550368 28350
rect 550048 28226 550368 28294
rect 550048 28170 550118 28226
rect 550174 28170 550242 28226
rect 550298 28170 550368 28226
rect 550048 28102 550368 28170
rect 550048 28046 550118 28102
rect 550174 28046 550242 28102
rect 550298 28046 550368 28102
rect 550048 27978 550368 28046
rect 550048 27922 550118 27978
rect 550174 27922 550242 27978
rect 550298 27922 550368 27978
rect 550048 27888 550368 27922
rect 585452 27972 585508 27982
rect 5418 22294 5514 22350
rect 5570 22294 5638 22350
rect 5694 22294 5762 22350
rect 5818 22294 5886 22350
rect 5942 22294 6038 22350
rect 5418 22226 6038 22294
rect 5418 22170 5514 22226
rect 5570 22170 5638 22226
rect 5694 22170 5762 22226
rect 5818 22170 5886 22226
rect 5942 22170 6038 22226
rect 5418 22102 6038 22170
rect 5418 22046 5514 22102
rect 5570 22046 5638 22102
rect 5694 22046 5762 22102
rect 5818 22046 5886 22102
rect 5942 22046 6038 22102
rect 5418 21978 6038 22046
rect 5418 21922 5514 21978
rect 5570 21922 5638 21978
rect 5694 21922 5762 21978
rect 5818 21922 5886 21978
rect 5942 21922 6038 21978
rect 5418 4350 6038 21922
rect 12448 22350 12768 22384
rect 12448 22294 12518 22350
rect 12574 22294 12642 22350
rect 12698 22294 12768 22350
rect 12448 22226 12768 22294
rect 12448 22170 12518 22226
rect 12574 22170 12642 22226
rect 12698 22170 12768 22226
rect 12448 22102 12768 22170
rect 12448 22046 12518 22102
rect 12574 22046 12642 22102
rect 12698 22046 12768 22102
rect 12448 21978 12768 22046
rect 12448 21922 12518 21978
rect 12574 21922 12642 21978
rect 12698 21922 12768 21978
rect 12448 21888 12768 21922
rect 43168 22350 43488 22384
rect 43168 22294 43238 22350
rect 43294 22294 43362 22350
rect 43418 22294 43488 22350
rect 43168 22226 43488 22294
rect 43168 22170 43238 22226
rect 43294 22170 43362 22226
rect 43418 22170 43488 22226
rect 43168 22102 43488 22170
rect 43168 22046 43238 22102
rect 43294 22046 43362 22102
rect 43418 22046 43488 22102
rect 43168 21978 43488 22046
rect 43168 21922 43238 21978
rect 43294 21922 43362 21978
rect 43418 21922 43488 21978
rect 43168 21888 43488 21922
rect 73888 22350 74208 22384
rect 73888 22294 73958 22350
rect 74014 22294 74082 22350
rect 74138 22294 74208 22350
rect 73888 22226 74208 22294
rect 73888 22170 73958 22226
rect 74014 22170 74082 22226
rect 74138 22170 74208 22226
rect 73888 22102 74208 22170
rect 73888 22046 73958 22102
rect 74014 22046 74082 22102
rect 74138 22046 74208 22102
rect 73888 21978 74208 22046
rect 73888 21922 73958 21978
rect 74014 21922 74082 21978
rect 74138 21922 74208 21978
rect 73888 21888 74208 21922
rect 104608 22350 104928 22384
rect 104608 22294 104678 22350
rect 104734 22294 104802 22350
rect 104858 22294 104928 22350
rect 104608 22226 104928 22294
rect 104608 22170 104678 22226
rect 104734 22170 104802 22226
rect 104858 22170 104928 22226
rect 104608 22102 104928 22170
rect 104608 22046 104678 22102
rect 104734 22046 104802 22102
rect 104858 22046 104928 22102
rect 104608 21978 104928 22046
rect 104608 21922 104678 21978
rect 104734 21922 104802 21978
rect 104858 21922 104928 21978
rect 104608 21888 104928 21922
rect 135328 22350 135648 22384
rect 135328 22294 135398 22350
rect 135454 22294 135522 22350
rect 135578 22294 135648 22350
rect 135328 22226 135648 22294
rect 135328 22170 135398 22226
rect 135454 22170 135522 22226
rect 135578 22170 135648 22226
rect 135328 22102 135648 22170
rect 135328 22046 135398 22102
rect 135454 22046 135522 22102
rect 135578 22046 135648 22102
rect 135328 21978 135648 22046
rect 135328 21922 135398 21978
rect 135454 21922 135522 21978
rect 135578 21922 135648 21978
rect 135328 21888 135648 21922
rect 166048 22350 166368 22384
rect 166048 22294 166118 22350
rect 166174 22294 166242 22350
rect 166298 22294 166368 22350
rect 166048 22226 166368 22294
rect 166048 22170 166118 22226
rect 166174 22170 166242 22226
rect 166298 22170 166368 22226
rect 166048 22102 166368 22170
rect 166048 22046 166118 22102
rect 166174 22046 166242 22102
rect 166298 22046 166368 22102
rect 166048 21978 166368 22046
rect 166048 21922 166118 21978
rect 166174 21922 166242 21978
rect 166298 21922 166368 21978
rect 166048 21888 166368 21922
rect 196768 22350 197088 22384
rect 196768 22294 196838 22350
rect 196894 22294 196962 22350
rect 197018 22294 197088 22350
rect 196768 22226 197088 22294
rect 196768 22170 196838 22226
rect 196894 22170 196962 22226
rect 197018 22170 197088 22226
rect 196768 22102 197088 22170
rect 196768 22046 196838 22102
rect 196894 22046 196962 22102
rect 197018 22046 197088 22102
rect 196768 21978 197088 22046
rect 196768 21922 196838 21978
rect 196894 21922 196962 21978
rect 197018 21922 197088 21978
rect 196768 21888 197088 21922
rect 227488 22350 227808 22384
rect 227488 22294 227558 22350
rect 227614 22294 227682 22350
rect 227738 22294 227808 22350
rect 227488 22226 227808 22294
rect 227488 22170 227558 22226
rect 227614 22170 227682 22226
rect 227738 22170 227808 22226
rect 227488 22102 227808 22170
rect 227488 22046 227558 22102
rect 227614 22046 227682 22102
rect 227738 22046 227808 22102
rect 227488 21978 227808 22046
rect 227488 21922 227558 21978
rect 227614 21922 227682 21978
rect 227738 21922 227808 21978
rect 227488 21888 227808 21922
rect 258208 22350 258528 22384
rect 258208 22294 258278 22350
rect 258334 22294 258402 22350
rect 258458 22294 258528 22350
rect 258208 22226 258528 22294
rect 258208 22170 258278 22226
rect 258334 22170 258402 22226
rect 258458 22170 258528 22226
rect 258208 22102 258528 22170
rect 258208 22046 258278 22102
rect 258334 22046 258402 22102
rect 258458 22046 258528 22102
rect 258208 21978 258528 22046
rect 258208 21922 258278 21978
rect 258334 21922 258402 21978
rect 258458 21922 258528 21978
rect 258208 21888 258528 21922
rect 288928 22350 289248 22384
rect 288928 22294 288998 22350
rect 289054 22294 289122 22350
rect 289178 22294 289248 22350
rect 288928 22226 289248 22294
rect 288928 22170 288998 22226
rect 289054 22170 289122 22226
rect 289178 22170 289248 22226
rect 288928 22102 289248 22170
rect 288928 22046 288998 22102
rect 289054 22046 289122 22102
rect 289178 22046 289248 22102
rect 288928 21978 289248 22046
rect 288928 21922 288998 21978
rect 289054 21922 289122 21978
rect 289178 21922 289248 21978
rect 288928 21888 289248 21922
rect 319648 22350 319968 22384
rect 319648 22294 319718 22350
rect 319774 22294 319842 22350
rect 319898 22294 319968 22350
rect 319648 22226 319968 22294
rect 319648 22170 319718 22226
rect 319774 22170 319842 22226
rect 319898 22170 319968 22226
rect 319648 22102 319968 22170
rect 319648 22046 319718 22102
rect 319774 22046 319842 22102
rect 319898 22046 319968 22102
rect 319648 21978 319968 22046
rect 319648 21922 319718 21978
rect 319774 21922 319842 21978
rect 319898 21922 319968 21978
rect 319648 21888 319968 21922
rect 350368 22350 350688 22384
rect 350368 22294 350438 22350
rect 350494 22294 350562 22350
rect 350618 22294 350688 22350
rect 350368 22226 350688 22294
rect 350368 22170 350438 22226
rect 350494 22170 350562 22226
rect 350618 22170 350688 22226
rect 350368 22102 350688 22170
rect 350368 22046 350438 22102
rect 350494 22046 350562 22102
rect 350618 22046 350688 22102
rect 350368 21978 350688 22046
rect 350368 21922 350438 21978
rect 350494 21922 350562 21978
rect 350618 21922 350688 21978
rect 350368 21888 350688 21922
rect 381088 22350 381408 22384
rect 381088 22294 381158 22350
rect 381214 22294 381282 22350
rect 381338 22294 381408 22350
rect 381088 22226 381408 22294
rect 381088 22170 381158 22226
rect 381214 22170 381282 22226
rect 381338 22170 381408 22226
rect 381088 22102 381408 22170
rect 381088 22046 381158 22102
rect 381214 22046 381282 22102
rect 381338 22046 381408 22102
rect 381088 21978 381408 22046
rect 381088 21922 381158 21978
rect 381214 21922 381282 21978
rect 381338 21922 381408 21978
rect 381088 21888 381408 21922
rect 411808 22350 412128 22384
rect 411808 22294 411878 22350
rect 411934 22294 412002 22350
rect 412058 22294 412128 22350
rect 411808 22226 412128 22294
rect 411808 22170 411878 22226
rect 411934 22170 412002 22226
rect 412058 22170 412128 22226
rect 411808 22102 412128 22170
rect 411808 22046 411878 22102
rect 411934 22046 412002 22102
rect 412058 22046 412128 22102
rect 411808 21978 412128 22046
rect 411808 21922 411878 21978
rect 411934 21922 412002 21978
rect 412058 21922 412128 21978
rect 411808 21888 412128 21922
rect 442528 22350 442848 22384
rect 442528 22294 442598 22350
rect 442654 22294 442722 22350
rect 442778 22294 442848 22350
rect 442528 22226 442848 22294
rect 442528 22170 442598 22226
rect 442654 22170 442722 22226
rect 442778 22170 442848 22226
rect 442528 22102 442848 22170
rect 442528 22046 442598 22102
rect 442654 22046 442722 22102
rect 442778 22046 442848 22102
rect 442528 21978 442848 22046
rect 442528 21922 442598 21978
rect 442654 21922 442722 21978
rect 442778 21922 442848 21978
rect 442528 21888 442848 21922
rect 473248 22350 473568 22384
rect 473248 22294 473318 22350
rect 473374 22294 473442 22350
rect 473498 22294 473568 22350
rect 473248 22226 473568 22294
rect 473248 22170 473318 22226
rect 473374 22170 473442 22226
rect 473498 22170 473568 22226
rect 473248 22102 473568 22170
rect 473248 22046 473318 22102
rect 473374 22046 473442 22102
rect 473498 22046 473568 22102
rect 473248 21978 473568 22046
rect 473248 21922 473318 21978
rect 473374 21922 473442 21978
rect 473498 21922 473568 21978
rect 473248 21888 473568 21922
rect 503968 22350 504288 22384
rect 503968 22294 504038 22350
rect 504094 22294 504162 22350
rect 504218 22294 504288 22350
rect 503968 22226 504288 22294
rect 503968 22170 504038 22226
rect 504094 22170 504162 22226
rect 504218 22170 504288 22226
rect 503968 22102 504288 22170
rect 503968 22046 504038 22102
rect 504094 22046 504162 22102
rect 504218 22046 504288 22102
rect 503968 21978 504288 22046
rect 503968 21922 504038 21978
rect 504094 21922 504162 21978
rect 504218 21922 504288 21978
rect 503968 21888 504288 21922
rect 534688 22350 535008 22384
rect 534688 22294 534758 22350
rect 534814 22294 534882 22350
rect 534938 22294 535008 22350
rect 534688 22226 535008 22294
rect 534688 22170 534758 22226
rect 534814 22170 534882 22226
rect 534938 22170 535008 22226
rect 534688 22102 535008 22170
rect 534688 22046 534758 22102
rect 534814 22046 534882 22102
rect 534938 22046 535008 22102
rect 534688 21978 535008 22046
rect 534688 21922 534758 21978
rect 534814 21922 534882 21978
rect 534938 21922 535008 21978
rect 534688 21888 535008 21922
rect 565408 22350 565728 22384
rect 565408 22294 565478 22350
rect 565534 22294 565602 22350
rect 565658 22294 565728 22350
rect 565408 22226 565728 22294
rect 565408 22170 565478 22226
rect 565534 22170 565602 22226
rect 565658 22170 565728 22226
rect 565408 22102 565728 22170
rect 565408 22046 565478 22102
rect 565534 22046 565602 22102
rect 565658 22046 565728 22102
rect 565408 21978 565728 22046
rect 565408 21922 565478 21978
rect 565534 21922 565602 21978
rect 565658 21922 565728 21978
rect 565408 21888 565728 21922
rect 585452 20356 585508 27916
rect 585452 20290 585508 20300
rect 589098 22350 589718 39922
rect 589098 22294 589194 22350
rect 589250 22294 589318 22350
rect 589374 22294 589442 22350
rect 589498 22294 589566 22350
rect 589622 22294 589718 22350
rect 589098 22226 589718 22294
rect 589098 22170 589194 22226
rect 589250 22170 589318 22226
rect 589374 22170 589442 22226
rect 589498 22170 589566 22226
rect 589622 22170 589718 22226
rect 589098 22102 589718 22170
rect 589098 22046 589194 22102
rect 589250 22046 589318 22102
rect 589374 22046 589442 22102
rect 589498 22046 589566 22102
rect 589622 22046 589718 22102
rect 589098 21978 589718 22046
rect 589098 21922 589194 21978
rect 589250 21922 589318 21978
rect 589374 21922 589442 21978
rect 589498 21922 589566 21978
rect 589622 21922 589718 21978
rect 6188 17668 6244 17678
rect 6188 8820 6244 17612
rect 6188 8754 6244 8764
rect 585452 17220 585508 17230
rect 5418 4294 5514 4350
rect 5570 4294 5638 4350
rect 5694 4294 5762 4350
rect 5818 4294 5886 4350
rect 5942 4294 6038 4350
rect 5418 4226 6038 4294
rect 5418 4170 5514 4226
rect 5570 4170 5638 4226
rect 5694 4170 5762 4226
rect 5818 4170 5886 4226
rect 5942 4170 6038 4226
rect 5418 4102 6038 4170
rect 5418 4046 5514 4102
rect 5570 4046 5638 4102
rect 5694 4046 5762 4102
rect 5818 4046 5886 4102
rect 5942 4046 6038 4102
rect 5418 3978 6038 4046
rect 5418 3922 5514 3978
rect 5570 3922 5638 3978
rect 5694 3922 5762 3978
rect 5818 3922 5886 3978
rect 5942 3922 6038 3978
rect 5418 -160 6038 3922
rect 5418 -216 5514 -160
rect 5570 -216 5638 -160
rect 5694 -216 5762 -160
rect 5818 -216 5886 -160
rect 5942 -216 6038 -160
rect 5418 -284 6038 -216
rect 5418 -340 5514 -284
rect 5570 -340 5638 -284
rect 5694 -340 5762 -284
rect 5818 -340 5886 -284
rect 5942 -340 6038 -284
rect 5418 -408 6038 -340
rect 5418 -464 5514 -408
rect 5570 -464 5638 -408
rect 5694 -464 5762 -408
rect 5818 -464 5886 -408
rect 5942 -464 6038 -408
rect 5418 -532 6038 -464
rect 5418 -588 5514 -532
rect 5570 -588 5638 -532
rect 5694 -588 5762 -532
rect 5818 -588 5886 -532
rect 5942 -588 6038 -532
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 -1296 -1120
rect -1916 -1244 -1296 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 -1296 -1244
rect -1916 -1368 -1296 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 -1296 -1368
rect -1916 -1492 -1296 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 -1296 -1492
rect -1916 -1644 -1296 -1548
rect 5418 -1644 6038 -588
rect 36138 4350 36758 7250
rect 36138 4294 36234 4350
rect 36290 4294 36358 4350
rect 36414 4294 36482 4350
rect 36538 4294 36606 4350
rect 36662 4294 36758 4350
rect 36138 4226 36758 4294
rect 36138 4170 36234 4226
rect 36290 4170 36358 4226
rect 36414 4170 36482 4226
rect 36538 4170 36606 4226
rect 36662 4170 36758 4226
rect 36138 4102 36758 4170
rect 36138 4046 36234 4102
rect 36290 4046 36358 4102
rect 36414 4046 36482 4102
rect 36538 4046 36606 4102
rect 36662 4046 36758 4102
rect 36138 3978 36758 4046
rect 36138 3922 36234 3978
rect 36290 3922 36358 3978
rect 36414 3922 36482 3978
rect 36538 3922 36606 3978
rect 36662 3922 36758 3978
rect 36138 -160 36758 3922
rect 36138 -216 36234 -160
rect 36290 -216 36358 -160
rect 36414 -216 36482 -160
rect 36538 -216 36606 -160
rect 36662 -216 36758 -160
rect 36138 -284 36758 -216
rect 36138 -340 36234 -284
rect 36290 -340 36358 -284
rect 36414 -340 36482 -284
rect 36538 -340 36606 -284
rect 36662 -340 36758 -284
rect 36138 -408 36758 -340
rect 36138 -464 36234 -408
rect 36290 -464 36358 -408
rect 36414 -464 36482 -408
rect 36538 -464 36606 -408
rect 36662 -464 36758 -408
rect 36138 -532 36758 -464
rect 36138 -588 36234 -532
rect 36290 -588 36358 -532
rect 36414 -588 36482 -532
rect 36538 -588 36606 -532
rect 36662 -588 36758 -532
rect 36138 -1644 36758 -588
rect 66858 4350 67478 7250
rect 66858 4294 66954 4350
rect 67010 4294 67078 4350
rect 67134 4294 67202 4350
rect 67258 4294 67326 4350
rect 67382 4294 67478 4350
rect 66858 4226 67478 4294
rect 66858 4170 66954 4226
rect 67010 4170 67078 4226
rect 67134 4170 67202 4226
rect 67258 4170 67326 4226
rect 67382 4170 67478 4226
rect 66858 4102 67478 4170
rect 66858 4046 66954 4102
rect 67010 4046 67078 4102
rect 67134 4046 67202 4102
rect 67258 4046 67326 4102
rect 67382 4046 67478 4102
rect 66858 3978 67478 4046
rect 66858 3922 66954 3978
rect 67010 3922 67078 3978
rect 67134 3922 67202 3978
rect 67258 3922 67326 3978
rect 67382 3922 67478 3978
rect 66858 -160 67478 3922
rect 66858 -216 66954 -160
rect 67010 -216 67078 -160
rect 67134 -216 67202 -160
rect 67258 -216 67326 -160
rect 67382 -216 67478 -160
rect 66858 -284 67478 -216
rect 66858 -340 66954 -284
rect 67010 -340 67078 -284
rect 67134 -340 67202 -284
rect 67258 -340 67326 -284
rect 67382 -340 67478 -284
rect 66858 -408 67478 -340
rect 66858 -464 66954 -408
rect 67010 -464 67078 -408
rect 67134 -464 67202 -408
rect 67258 -464 67326 -408
rect 67382 -464 67478 -408
rect 66858 -532 67478 -464
rect 66858 -588 66954 -532
rect 67010 -588 67078 -532
rect 67134 -588 67202 -532
rect 67258 -588 67326 -532
rect 67382 -588 67478 -532
rect 66858 -1644 67478 -588
rect 97578 4350 98198 7250
rect 97578 4294 97674 4350
rect 97730 4294 97798 4350
rect 97854 4294 97922 4350
rect 97978 4294 98046 4350
rect 98102 4294 98198 4350
rect 97578 4226 98198 4294
rect 97578 4170 97674 4226
rect 97730 4170 97798 4226
rect 97854 4170 97922 4226
rect 97978 4170 98046 4226
rect 98102 4170 98198 4226
rect 97578 4102 98198 4170
rect 97578 4046 97674 4102
rect 97730 4046 97798 4102
rect 97854 4046 97922 4102
rect 97978 4046 98046 4102
rect 98102 4046 98198 4102
rect 97578 3978 98198 4046
rect 97578 3922 97674 3978
rect 97730 3922 97798 3978
rect 97854 3922 97922 3978
rect 97978 3922 98046 3978
rect 98102 3922 98198 3978
rect 97578 -160 98198 3922
rect 97578 -216 97674 -160
rect 97730 -216 97798 -160
rect 97854 -216 97922 -160
rect 97978 -216 98046 -160
rect 98102 -216 98198 -160
rect 97578 -284 98198 -216
rect 97578 -340 97674 -284
rect 97730 -340 97798 -284
rect 97854 -340 97922 -284
rect 97978 -340 98046 -284
rect 98102 -340 98198 -284
rect 97578 -408 98198 -340
rect 97578 -464 97674 -408
rect 97730 -464 97798 -408
rect 97854 -464 97922 -408
rect 97978 -464 98046 -408
rect 98102 -464 98198 -408
rect 97578 -532 98198 -464
rect 97578 -588 97674 -532
rect 97730 -588 97798 -532
rect 97854 -588 97922 -532
rect 97978 -588 98046 -532
rect 98102 -588 98198 -532
rect 97578 -1644 98198 -588
rect 128298 4350 128918 7250
rect 128298 4294 128394 4350
rect 128450 4294 128518 4350
rect 128574 4294 128642 4350
rect 128698 4294 128766 4350
rect 128822 4294 128918 4350
rect 128298 4226 128918 4294
rect 128298 4170 128394 4226
rect 128450 4170 128518 4226
rect 128574 4170 128642 4226
rect 128698 4170 128766 4226
rect 128822 4170 128918 4226
rect 128298 4102 128918 4170
rect 128298 4046 128394 4102
rect 128450 4046 128518 4102
rect 128574 4046 128642 4102
rect 128698 4046 128766 4102
rect 128822 4046 128918 4102
rect 128298 3978 128918 4046
rect 128298 3922 128394 3978
rect 128450 3922 128518 3978
rect 128574 3922 128642 3978
rect 128698 3922 128766 3978
rect 128822 3922 128918 3978
rect 128298 -160 128918 3922
rect 128298 -216 128394 -160
rect 128450 -216 128518 -160
rect 128574 -216 128642 -160
rect 128698 -216 128766 -160
rect 128822 -216 128918 -160
rect 128298 -284 128918 -216
rect 128298 -340 128394 -284
rect 128450 -340 128518 -284
rect 128574 -340 128642 -284
rect 128698 -340 128766 -284
rect 128822 -340 128918 -284
rect 128298 -408 128918 -340
rect 128298 -464 128394 -408
rect 128450 -464 128518 -408
rect 128574 -464 128642 -408
rect 128698 -464 128766 -408
rect 128822 -464 128918 -408
rect 128298 -532 128918 -464
rect 128298 -588 128394 -532
rect 128450 -588 128518 -532
rect 128574 -588 128642 -532
rect 128698 -588 128766 -532
rect 128822 -588 128918 -532
rect 128298 -1644 128918 -588
rect 159018 4350 159638 7250
rect 159018 4294 159114 4350
rect 159170 4294 159238 4350
rect 159294 4294 159362 4350
rect 159418 4294 159486 4350
rect 159542 4294 159638 4350
rect 159018 4226 159638 4294
rect 159018 4170 159114 4226
rect 159170 4170 159238 4226
rect 159294 4170 159362 4226
rect 159418 4170 159486 4226
rect 159542 4170 159638 4226
rect 159018 4102 159638 4170
rect 159018 4046 159114 4102
rect 159170 4046 159238 4102
rect 159294 4046 159362 4102
rect 159418 4046 159486 4102
rect 159542 4046 159638 4102
rect 159018 3978 159638 4046
rect 159018 3922 159114 3978
rect 159170 3922 159238 3978
rect 159294 3922 159362 3978
rect 159418 3922 159486 3978
rect 159542 3922 159638 3978
rect 159018 -160 159638 3922
rect 159018 -216 159114 -160
rect 159170 -216 159238 -160
rect 159294 -216 159362 -160
rect 159418 -216 159486 -160
rect 159542 -216 159638 -160
rect 159018 -284 159638 -216
rect 159018 -340 159114 -284
rect 159170 -340 159238 -284
rect 159294 -340 159362 -284
rect 159418 -340 159486 -284
rect 159542 -340 159638 -284
rect 159018 -408 159638 -340
rect 159018 -464 159114 -408
rect 159170 -464 159238 -408
rect 159294 -464 159362 -408
rect 159418 -464 159486 -408
rect 159542 -464 159638 -408
rect 159018 -532 159638 -464
rect 159018 -588 159114 -532
rect 159170 -588 159238 -532
rect 159294 -588 159362 -532
rect 159418 -588 159486 -532
rect 159542 -588 159638 -532
rect 159018 -1644 159638 -588
rect 189738 4350 190358 7250
rect 189738 4294 189834 4350
rect 189890 4294 189958 4350
rect 190014 4294 190082 4350
rect 190138 4294 190206 4350
rect 190262 4294 190358 4350
rect 189738 4226 190358 4294
rect 189738 4170 189834 4226
rect 189890 4170 189958 4226
rect 190014 4170 190082 4226
rect 190138 4170 190206 4226
rect 190262 4170 190358 4226
rect 189738 4102 190358 4170
rect 189738 4046 189834 4102
rect 189890 4046 189958 4102
rect 190014 4046 190082 4102
rect 190138 4046 190206 4102
rect 190262 4046 190358 4102
rect 189738 3978 190358 4046
rect 189738 3922 189834 3978
rect 189890 3922 189958 3978
rect 190014 3922 190082 3978
rect 190138 3922 190206 3978
rect 190262 3922 190358 3978
rect 189738 -160 190358 3922
rect 189738 -216 189834 -160
rect 189890 -216 189958 -160
rect 190014 -216 190082 -160
rect 190138 -216 190206 -160
rect 190262 -216 190358 -160
rect 189738 -284 190358 -216
rect 189738 -340 189834 -284
rect 189890 -340 189958 -284
rect 190014 -340 190082 -284
rect 190138 -340 190206 -284
rect 190262 -340 190358 -284
rect 189738 -408 190358 -340
rect 189738 -464 189834 -408
rect 189890 -464 189958 -408
rect 190014 -464 190082 -408
rect 190138 -464 190206 -408
rect 190262 -464 190358 -408
rect 189738 -532 190358 -464
rect 189738 -588 189834 -532
rect 189890 -588 189958 -532
rect 190014 -588 190082 -532
rect 190138 -588 190206 -532
rect 190262 -588 190358 -532
rect 189738 -1644 190358 -588
rect 220458 4350 221078 7250
rect 220458 4294 220554 4350
rect 220610 4294 220678 4350
rect 220734 4294 220802 4350
rect 220858 4294 220926 4350
rect 220982 4294 221078 4350
rect 220458 4226 221078 4294
rect 220458 4170 220554 4226
rect 220610 4170 220678 4226
rect 220734 4170 220802 4226
rect 220858 4170 220926 4226
rect 220982 4170 221078 4226
rect 220458 4102 221078 4170
rect 220458 4046 220554 4102
rect 220610 4046 220678 4102
rect 220734 4046 220802 4102
rect 220858 4046 220926 4102
rect 220982 4046 221078 4102
rect 220458 3978 221078 4046
rect 220458 3922 220554 3978
rect 220610 3922 220678 3978
rect 220734 3922 220802 3978
rect 220858 3922 220926 3978
rect 220982 3922 221078 3978
rect 220458 -160 221078 3922
rect 220458 -216 220554 -160
rect 220610 -216 220678 -160
rect 220734 -216 220802 -160
rect 220858 -216 220926 -160
rect 220982 -216 221078 -160
rect 220458 -284 221078 -216
rect 220458 -340 220554 -284
rect 220610 -340 220678 -284
rect 220734 -340 220802 -284
rect 220858 -340 220926 -284
rect 220982 -340 221078 -284
rect 220458 -408 221078 -340
rect 220458 -464 220554 -408
rect 220610 -464 220678 -408
rect 220734 -464 220802 -408
rect 220858 -464 220926 -408
rect 220982 -464 221078 -408
rect 220458 -532 221078 -464
rect 220458 -588 220554 -532
rect 220610 -588 220678 -532
rect 220734 -588 220802 -532
rect 220858 -588 220926 -532
rect 220982 -588 221078 -532
rect 220458 -1644 221078 -588
rect 251178 4350 251798 7250
rect 251178 4294 251274 4350
rect 251330 4294 251398 4350
rect 251454 4294 251522 4350
rect 251578 4294 251646 4350
rect 251702 4294 251798 4350
rect 251178 4226 251798 4294
rect 251178 4170 251274 4226
rect 251330 4170 251398 4226
rect 251454 4170 251522 4226
rect 251578 4170 251646 4226
rect 251702 4170 251798 4226
rect 251178 4102 251798 4170
rect 251178 4046 251274 4102
rect 251330 4046 251398 4102
rect 251454 4046 251522 4102
rect 251578 4046 251646 4102
rect 251702 4046 251798 4102
rect 251178 3978 251798 4046
rect 251178 3922 251274 3978
rect 251330 3922 251398 3978
rect 251454 3922 251522 3978
rect 251578 3922 251646 3978
rect 251702 3922 251798 3978
rect 251178 -160 251798 3922
rect 251178 -216 251274 -160
rect 251330 -216 251398 -160
rect 251454 -216 251522 -160
rect 251578 -216 251646 -160
rect 251702 -216 251798 -160
rect 251178 -284 251798 -216
rect 251178 -340 251274 -284
rect 251330 -340 251398 -284
rect 251454 -340 251522 -284
rect 251578 -340 251646 -284
rect 251702 -340 251798 -284
rect 251178 -408 251798 -340
rect 251178 -464 251274 -408
rect 251330 -464 251398 -408
rect 251454 -464 251522 -408
rect 251578 -464 251646 -408
rect 251702 -464 251798 -408
rect 251178 -532 251798 -464
rect 251178 -588 251274 -532
rect 251330 -588 251398 -532
rect 251454 -588 251522 -532
rect 251578 -588 251646 -532
rect 251702 -588 251798 -532
rect 251178 -1644 251798 -588
rect 281898 4350 282518 7250
rect 281898 4294 281994 4350
rect 282050 4294 282118 4350
rect 282174 4294 282242 4350
rect 282298 4294 282366 4350
rect 282422 4294 282518 4350
rect 281898 4226 282518 4294
rect 281898 4170 281994 4226
rect 282050 4170 282118 4226
rect 282174 4170 282242 4226
rect 282298 4170 282366 4226
rect 282422 4170 282518 4226
rect 281898 4102 282518 4170
rect 281898 4046 281994 4102
rect 282050 4046 282118 4102
rect 282174 4046 282242 4102
rect 282298 4046 282366 4102
rect 282422 4046 282518 4102
rect 281898 3978 282518 4046
rect 281898 3922 281994 3978
rect 282050 3922 282118 3978
rect 282174 3922 282242 3978
rect 282298 3922 282366 3978
rect 282422 3922 282518 3978
rect 281898 -160 282518 3922
rect 281898 -216 281994 -160
rect 282050 -216 282118 -160
rect 282174 -216 282242 -160
rect 282298 -216 282366 -160
rect 282422 -216 282518 -160
rect 281898 -284 282518 -216
rect 281898 -340 281994 -284
rect 282050 -340 282118 -284
rect 282174 -340 282242 -284
rect 282298 -340 282366 -284
rect 282422 -340 282518 -284
rect 281898 -408 282518 -340
rect 281898 -464 281994 -408
rect 282050 -464 282118 -408
rect 282174 -464 282242 -408
rect 282298 -464 282366 -408
rect 282422 -464 282518 -408
rect 281898 -532 282518 -464
rect 281898 -588 281994 -532
rect 282050 -588 282118 -532
rect 282174 -588 282242 -532
rect 282298 -588 282366 -532
rect 282422 -588 282518 -532
rect 281898 -1644 282518 -588
rect 312618 4350 313238 7250
rect 312618 4294 312714 4350
rect 312770 4294 312838 4350
rect 312894 4294 312962 4350
rect 313018 4294 313086 4350
rect 313142 4294 313238 4350
rect 312618 4226 313238 4294
rect 312618 4170 312714 4226
rect 312770 4170 312838 4226
rect 312894 4170 312962 4226
rect 313018 4170 313086 4226
rect 313142 4170 313238 4226
rect 312618 4102 313238 4170
rect 312618 4046 312714 4102
rect 312770 4046 312838 4102
rect 312894 4046 312962 4102
rect 313018 4046 313086 4102
rect 313142 4046 313238 4102
rect 312618 3978 313238 4046
rect 312618 3922 312714 3978
rect 312770 3922 312838 3978
rect 312894 3922 312962 3978
rect 313018 3922 313086 3978
rect 313142 3922 313238 3978
rect 312618 -160 313238 3922
rect 312618 -216 312714 -160
rect 312770 -216 312838 -160
rect 312894 -216 312962 -160
rect 313018 -216 313086 -160
rect 313142 -216 313238 -160
rect 312618 -284 313238 -216
rect 312618 -340 312714 -284
rect 312770 -340 312838 -284
rect 312894 -340 312962 -284
rect 313018 -340 313086 -284
rect 313142 -340 313238 -284
rect 312618 -408 313238 -340
rect 312618 -464 312714 -408
rect 312770 -464 312838 -408
rect 312894 -464 312962 -408
rect 313018 -464 313086 -408
rect 313142 -464 313238 -408
rect 312618 -532 313238 -464
rect 312618 -588 312714 -532
rect 312770 -588 312838 -532
rect 312894 -588 312962 -532
rect 313018 -588 313086 -532
rect 313142 -588 313238 -532
rect 312618 -1644 313238 -588
rect 343338 4350 343958 7250
rect 343338 4294 343434 4350
rect 343490 4294 343558 4350
rect 343614 4294 343682 4350
rect 343738 4294 343806 4350
rect 343862 4294 343958 4350
rect 343338 4226 343958 4294
rect 343338 4170 343434 4226
rect 343490 4170 343558 4226
rect 343614 4170 343682 4226
rect 343738 4170 343806 4226
rect 343862 4170 343958 4226
rect 343338 4102 343958 4170
rect 343338 4046 343434 4102
rect 343490 4046 343558 4102
rect 343614 4046 343682 4102
rect 343738 4046 343806 4102
rect 343862 4046 343958 4102
rect 343338 3978 343958 4046
rect 343338 3922 343434 3978
rect 343490 3922 343558 3978
rect 343614 3922 343682 3978
rect 343738 3922 343806 3978
rect 343862 3922 343958 3978
rect 343338 -160 343958 3922
rect 343338 -216 343434 -160
rect 343490 -216 343558 -160
rect 343614 -216 343682 -160
rect 343738 -216 343806 -160
rect 343862 -216 343958 -160
rect 343338 -284 343958 -216
rect 343338 -340 343434 -284
rect 343490 -340 343558 -284
rect 343614 -340 343682 -284
rect 343738 -340 343806 -284
rect 343862 -340 343958 -284
rect 343338 -408 343958 -340
rect 343338 -464 343434 -408
rect 343490 -464 343558 -408
rect 343614 -464 343682 -408
rect 343738 -464 343806 -408
rect 343862 -464 343958 -408
rect 343338 -532 343958 -464
rect 343338 -588 343434 -532
rect 343490 -588 343558 -532
rect 343614 -588 343682 -532
rect 343738 -588 343806 -532
rect 343862 -588 343958 -532
rect 343338 -1644 343958 -588
rect 374058 4350 374678 7250
rect 374058 4294 374154 4350
rect 374210 4294 374278 4350
rect 374334 4294 374402 4350
rect 374458 4294 374526 4350
rect 374582 4294 374678 4350
rect 374058 4226 374678 4294
rect 374058 4170 374154 4226
rect 374210 4170 374278 4226
rect 374334 4170 374402 4226
rect 374458 4170 374526 4226
rect 374582 4170 374678 4226
rect 374058 4102 374678 4170
rect 374058 4046 374154 4102
rect 374210 4046 374278 4102
rect 374334 4046 374402 4102
rect 374458 4046 374526 4102
rect 374582 4046 374678 4102
rect 374058 3978 374678 4046
rect 374058 3922 374154 3978
rect 374210 3922 374278 3978
rect 374334 3922 374402 3978
rect 374458 3922 374526 3978
rect 374582 3922 374678 3978
rect 374058 -160 374678 3922
rect 374058 -216 374154 -160
rect 374210 -216 374278 -160
rect 374334 -216 374402 -160
rect 374458 -216 374526 -160
rect 374582 -216 374678 -160
rect 374058 -284 374678 -216
rect 374058 -340 374154 -284
rect 374210 -340 374278 -284
rect 374334 -340 374402 -284
rect 374458 -340 374526 -284
rect 374582 -340 374678 -284
rect 374058 -408 374678 -340
rect 374058 -464 374154 -408
rect 374210 -464 374278 -408
rect 374334 -464 374402 -408
rect 374458 -464 374526 -408
rect 374582 -464 374678 -408
rect 374058 -532 374678 -464
rect 374058 -588 374154 -532
rect 374210 -588 374278 -532
rect 374334 -588 374402 -532
rect 374458 -588 374526 -532
rect 374582 -588 374678 -532
rect 374058 -1644 374678 -588
rect 404778 4350 405398 7250
rect 404778 4294 404874 4350
rect 404930 4294 404998 4350
rect 405054 4294 405122 4350
rect 405178 4294 405246 4350
rect 405302 4294 405398 4350
rect 404778 4226 405398 4294
rect 404778 4170 404874 4226
rect 404930 4170 404998 4226
rect 405054 4170 405122 4226
rect 405178 4170 405246 4226
rect 405302 4170 405398 4226
rect 404778 4102 405398 4170
rect 404778 4046 404874 4102
rect 404930 4046 404998 4102
rect 405054 4046 405122 4102
rect 405178 4046 405246 4102
rect 405302 4046 405398 4102
rect 404778 3978 405398 4046
rect 404778 3922 404874 3978
rect 404930 3922 404998 3978
rect 405054 3922 405122 3978
rect 405178 3922 405246 3978
rect 405302 3922 405398 3978
rect 404778 -160 405398 3922
rect 404778 -216 404874 -160
rect 404930 -216 404998 -160
rect 405054 -216 405122 -160
rect 405178 -216 405246 -160
rect 405302 -216 405398 -160
rect 404778 -284 405398 -216
rect 404778 -340 404874 -284
rect 404930 -340 404998 -284
rect 405054 -340 405122 -284
rect 405178 -340 405246 -284
rect 405302 -340 405398 -284
rect 404778 -408 405398 -340
rect 404778 -464 404874 -408
rect 404930 -464 404998 -408
rect 405054 -464 405122 -408
rect 405178 -464 405246 -408
rect 405302 -464 405398 -408
rect 404778 -532 405398 -464
rect 404778 -588 404874 -532
rect 404930 -588 404998 -532
rect 405054 -588 405122 -532
rect 405178 -588 405246 -532
rect 405302 -588 405398 -532
rect 404778 -1644 405398 -588
rect 435498 4350 436118 7250
rect 435498 4294 435594 4350
rect 435650 4294 435718 4350
rect 435774 4294 435842 4350
rect 435898 4294 435966 4350
rect 436022 4294 436118 4350
rect 435498 4226 436118 4294
rect 435498 4170 435594 4226
rect 435650 4170 435718 4226
rect 435774 4170 435842 4226
rect 435898 4170 435966 4226
rect 436022 4170 436118 4226
rect 435498 4102 436118 4170
rect 435498 4046 435594 4102
rect 435650 4046 435718 4102
rect 435774 4046 435842 4102
rect 435898 4046 435966 4102
rect 436022 4046 436118 4102
rect 435498 3978 436118 4046
rect 435498 3922 435594 3978
rect 435650 3922 435718 3978
rect 435774 3922 435842 3978
rect 435898 3922 435966 3978
rect 436022 3922 436118 3978
rect 435498 -160 436118 3922
rect 435498 -216 435594 -160
rect 435650 -216 435718 -160
rect 435774 -216 435842 -160
rect 435898 -216 435966 -160
rect 436022 -216 436118 -160
rect 435498 -284 436118 -216
rect 435498 -340 435594 -284
rect 435650 -340 435718 -284
rect 435774 -340 435842 -284
rect 435898 -340 435966 -284
rect 436022 -340 436118 -284
rect 435498 -408 436118 -340
rect 435498 -464 435594 -408
rect 435650 -464 435718 -408
rect 435774 -464 435842 -408
rect 435898 -464 435966 -408
rect 436022 -464 436118 -408
rect 435498 -532 436118 -464
rect 435498 -588 435594 -532
rect 435650 -588 435718 -532
rect 435774 -588 435842 -532
rect 435898 -588 435966 -532
rect 436022 -588 436118 -532
rect 435498 -1644 436118 -588
rect 466218 4350 466838 7250
rect 466218 4294 466314 4350
rect 466370 4294 466438 4350
rect 466494 4294 466562 4350
rect 466618 4294 466686 4350
rect 466742 4294 466838 4350
rect 466218 4226 466838 4294
rect 466218 4170 466314 4226
rect 466370 4170 466438 4226
rect 466494 4170 466562 4226
rect 466618 4170 466686 4226
rect 466742 4170 466838 4226
rect 466218 4102 466838 4170
rect 466218 4046 466314 4102
rect 466370 4046 466438 4102
rect 466494 4046 466562 4102
rect 466618 4046 466686 4102
rect 466742 4046 466838 4102
rect 466218 3978 466838 4046
rect 466218 3922 466314 3978
rect 466370 3922 466438 3978
rect 466494 3922 466562 3978
rect 466618 3922 466686 3978
rect 466742 3922 466838 3978
rect 466218 -160 466838 3922
rect 466218 -216 466314 -160
rect 466370 -216 466438 -160
rect 466494 -216 466562 -160
rect 466618 -216 466686 -160
rect 466742 -216 466838 -160
rect 466218 -284 466838 -216
rect 466218 -340 466314 -284
rect 466370 -340 466438 -284
rect 466494 -340 466562 -284
rect 466618 -340 466686 -284
rect 466742 -340 466838 -284
rect 466218 -408 466838 -340
rect 466218 -464 466314 -408
rect 466370 -464 466438 -408
rect 466494 -464 466562 -408
rect 466618 -464 466686 -408
rect 466742 -464 466838 -408
rect 466218 -532 466838 -464
rect 466218 -588 466314 -532
rect 466370 -588 466438 -532
rect 466494 -588 466562 -532
rect 466618 -588 466686 -532
rect 466742 -588 466838 -532
rect 466218 -1644 466838 -588
rect 496938 4350 497558 7250
rect 496938 4294 497034 4350
rect 497090 4294 497158 4350
rect 497214 4294 497282 4350
rect 497338 4294 497406 4350
rect 497462 4294 497558 4350
rect 496938 4226 497558 4294
rect 496938 4170 497034 4226
rect 497090 4170 497158 4226
rect 497214 4170 497282 4226
rect 497338 4170 497406 4226
rect 497462 4170 497558 4226
rect 496938 4102 497558 4170
rect 496938 4046 497034 4102
rect 497090 4046 497158 4102
rect 497214 4046 497282 4102
rect 497338 4046 497406 4102
rect 497462 4046 497558 4102
rect 496938 3978 497558 4046
rect 496938 3922 497034 3978
rect 497090 3922 497158 3978
rect 497214 3922 497282 3978
rect 497338 3922 497406 3978
rect 497462 3922 497558 3978
rect 496938 -160 497558 3922
rect 496938 -216 497034 -160
rect 497090 -216 497158 -160
rect 497214 -216 497282 -160
rect 497338 -216 497406 -160
rect 497462 -216 497558 -160
rect 496938 -284 497558 -216
rect 496938 -340 497034 -284
rect 497090 -340 497158 -284
rect 497214 -340 497282 -284
rect 497338 -340 497406 -284
rect 497462 -340 497558 -284
rect 496938 -408 497558 -340
rect 496938 -464 497034 -408
rect 497090 -464 497158 -408
rect 497214 -464 497282 -408
rect 497338 -464 497406 -408
rect 497462 -464 497558 -408
rect 496938 -532 497558 -464
rect 496938 -588 497034 -532
rect 497090 -588 497158 -532
rect 497214 -588 497282 -532
rect 497338 -588 497406 -532
rect 497462 -588 497558 -532
rect 496938 -1644 497558 -588
rect 527658 4350 528278 7250
rect 557452 6580 557508 6590
rect 557452 4978 557508 6524
rect 557452 4912 557508 4922
rect 527658 4294 527754 4350
rect 527810 4294 527878 4350
rect 527934 4294 528002 4350
rect 528058 4294 528126 4350
rect 528182 4294 528278 4350
rect 527658 4226 528278 4294
rect 527658 4170 527754 4226
rect 527810 4170 527878 4226
rect 527934 4170 528002 4226
rect 528058 4170 528126 4226
rect 528182 4170 528278 4226
rect 527658 4102 528278 4170
rect 527658 4046 527754 4102
rect 527810 4046 527878 4102
rect 527934 4046 528002 4102
rect 528058 4046 528126 4102
rect 528182 4046 528278 4102
rect 527658 3978 528278 4046
rect 527658 3922 527754 3978
rect 527810 3922 527878 3978
rect 527934 3922 528002 3978
rect 528058 3922 528126 3978
rect 528182 3922 528278 3978
rect 527658 -160 528278 3922
rect 527658 -216 527754 -160
rect 527810 -216 527878 -160
rect 527934 -216 528002 -160
rect 528058 -216 528126 -160
rect 528182 -216 528278 -160
rect 527658 -284 528278 -216
rect 527658 -340 527754 -284
rect 527810 -340 527878 -284
rect 527934 -340 528002 -284
rect 528058 -340 528126 -284
rect 528182 -340 528278 -284
rect 527658 -408 528278 -340
rect 527658 -464 527754 -408
rect 527810 -464 527878 -408
rect 527934 -464 528002 -408
rect 528058 -464 528126 -408
rect 528182 -464 528278 -408
rect 527658 -532 528278 -464
rect 527658 -588 527754 -532
rect 527810 -588 527878 -532
rect 527934 -588 528002 -532
rect 528058 -588 528126 -532
rect 528182 -588 528278 -532
rect 527658 -1644 528278 -588
rect 558378 4350 558998 7250
rect 585452 7140 585508 17164
rect 585452 7074 585508 7084
rect 561036 6468 561092 6478
rect 561036 4798 561092 6412
rect 561036 4732 561092 4742
rect 576828 4978 576884 4988
rect 558378 4294 558474 4350
rect 558530 4294 558598 4350
rect 558654 4294 558722 4350
rect 558778 4294 558846 4350
rect 558902 4294 558998 4350
rect 558378 4226 558998 4294
rect 558378 4170 558474 4226
rect 558530 4170 558598 4226
rect 558654 4170 558722 4226
rect 558778 4170 558846 4226
rect 558902 4170 558998 4226
rect 558378 4102 558998 4170
rect 558378 4046 558474 4102
rect 558530 4046 558598 4102
rect 558654 4046 558722 4102
rect 558778 4046 558846 4102
rect 558902 4046 558998 4102
rect 558378 3978 558998 4046
rect 558378 3922 558474 3978
rect 558530 3922 558598 3978
rect 558654 3922 558722 3978
rect 558778 3922 558846 3978
rect 558902 3922 558998 3978
rect 558378 -160 558998 3922
rect 576828 3444 576884 4922
rect 576828 3378 576884 3388
rect 580636 4798 580692 4808
rect 580636 3444 580692 4742
rect 580636 3378 580692 3388
rect 589098 4350 589718 21922
rect 589098 4294 589194 4350
rect 589250 4294 589318 4350
rect 589374 4294 589442 4350
rect 589498 4294 589566 4350
rect 589622 4294 589718 4350
rect 589098 4226 589718 4294
rect 589098 4170 589194 4226
rect 589250 4170 589318 4226
rect 589374 4170 589442 4226
rect 589498 4170 589566 4226
rect 589622 4170 589718 4226
rect 589098 4102 589718 4170
rect 589098 4046 589194 4102
rect 589250 4046 589318 4102
rect 589374 4046 589442 4102
rect 589498 4046 589566 4102
rect 589622 4046 589718 4102
rect 589098 3978 589718 4046
rect 589098 3922 589194 3978
rect 589250 3922 589318 3978
rect 589374 3922 589442 3978
rect 589498 3922 589566 3978
rect 589622 3922 589718 3978
rect 558378 -216 558474 -160
rect 558530 -216 558598 -160
rect 558654 -216 558722 -160
rect 558778 -216 558846 -160
rect 558902 -216 558998 -160
rect 558378 -284 558998 -216
rect 558378 -340 558474 -284
rect 558530 -340 558598 -284
rect 558654 -340 558722 -284
rect 558778 -340 558846 -284
rect 558902 -340 558998 -284
rect 558378 -408 558998 -340
rect 558378 -464 558474 -408
rect 558530 -464 558598 -408
rect 558654 -464 558722 -408
rect 558778 -464 558846 -408
rect 558902 -464 558998 -408
rect 558378 -532 558998 -464
rect 558378 -588 558474 -532
rect 558530 -588 558598 -532
rect 558654 -588 558722 -532
rect 558778 -588 558846 -532
rect 558902 -588 558998 -532
rect 558378 -1644 558998 -588
rect 589098 -160 589718 3922
rect 589098 -216 589194 -160
rect 589250 -216 589318 -160
rect 589374 -216 589442 -160
rect 589498 -216 589566 -160
rect 589622 -216 589718 -160
rect 589098 -284 589718 -216
rect 589098 -340 589194 -284
rect 589250 -340 589318 -284
rect 589374 -340 589442 -284
rect 589498 -340 589566 -284
rect 589622 -340 589718 -284
rect 589098 -408 589718 -340
rect 589098 -464 589194 -408
rect 589250 -464 589318 -408
rect 589374 -464 589442 -408
rect 589498 -464 589566 -408
rect 589622 -464 589718 -408
rect 589098 -532 589718 -464
rect 589098 -588 589194 -532
rect 589250 -588 589318 -532
rect 589374 -588 589442 -532
rect 589498 -588 589566 -532
rect 589622 -588 589718 -532
rect 589098 -1644 589718 -588
rect 592818 46350 593438 63922
rect 592818 46294 592914 46350
rect 592970 46294 593038 46350
rect 593094 46294 593162 46350
rect 593218 46294 593286 46350
rect 593342 46294 593438 46350
rect 592818 46226 593438 46294
rect 592818 46170 592914 46226
rect 592970 46170 593038 46226
rect 593094 46170 593162 46226
rect 593218 46170 593286 46226
rect 593342 46170 593438 46226
rect 592818 46102 593438 46170
rect 592818 46046 592914 46102
rect 592970 46046 593038 46102
rect 593094 46046 593162 46102
rect 593218 46046 593286 46102
rect 593342 46046 593438 46102
rect 592818 45978 593438 46046
rect 592818 45922 592914 45978
rect 592970 45922 593038 45978
rect 593094 45922 593162 45978
rect 593218 45922 593286 45978
rect 593342 45922 593438 45978
rect 592818 28350 593438 45922
rect 592818 28294 592914 28350
rect 592970 28294 593038 28350
rect 593094 28294 593162 28350
rect 593218 28294 593286 28350
rect 593342 28294 593438 28350
rect 592818 28226 593438 28294
rect 592818 28170 592914 28226
rect 592970 28170 593038 28226
rect 593094 28170 593162 28226
rect 593218 28170 593286 28226
rect 593342 28170 593438 28226
rect 592818 28102 593438 28170
rect 592818 28046 592914 28102
rect 592970 28046 593038 28102
rect 593094 28046 593162 28102
rect 593218 28046 593286 28102
rect 593342 28046 593438 28102
rect 592818 27978 593438 28046
rect 592818 27922 592914 27978
rect 592970 27922 593038 27978
rect 593094 27922 593162 27978
rect 593218 27922 593286 27978
rect 593342 27922 593438 27978
rect 592818 10350 593438 27922
rect 592818 10294 592914 10350
rect 592970 10294 593038 10350
rect 593094 10294 593162 10350
rect 593218 10294 593286 10350
rect 593342 10294 593438 10350
rect 592818 10226 593438 10294
rect 592818 10170 592914 10226
rect 592970 10170 593038 10226
rect 593094 10170 593162 10226
rect 593218 10170 593286 10226
rect 593342 10170 593438 10226
rect 592818 10102 593438 10170
rect 592818 10046 592914 10102
rect 592970 10046 593038 10102
rect 593094 10046 593162 10102
rect 593218 10046 593286 10102
rect 593342 10046 593438 10102
rect 592818 9978 593438 10046
rect 592818 9922 592914 9978
rect 592970 9922 593038 9978
rect 593094 9922 593162 9978
rect 593218 9922 593286 9978
rect 593342 9922 593438 9978
rect 592818 -1120 593438 9922
rect 596400 597212 597020 597308
rect 596400 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect 596400 597088 597020 597156
rect 596400 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect 596400 596964 597020 597032
rect 596400 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect 596400 596840 597020 596908
rect 596400 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect 596400 580350 597020 596784
rect 596400 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597020 580350
rect 596400 580226 597020 580294
rect 596400 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597020 580226
rect 596400 580102 597020 580170
rect 596400 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597020 580102
rect 596400 579978 597020 580046
rect 596400 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597020 579978
rect 596400 562350 597020 579922
rect 596400 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597020 562350
rect 596400 562226 597020 562294
rect 596400 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597020 562226
rect 596400 562102 597020 562170
rect 596400 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597020 562102
rect 596400 561978 597020 562046
rect 596400 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597020 561978
rect 596400 544350 597020 561922
rect 596400 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597020 544350
rect 596400 544226 597020 544294
rect 596400 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597020 544226
rect 596400 544102 597020 544170
rect 596400 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597020 544102
rect 596400 543978 597020 544046
rect 596400 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597020 543978
rect 596400 526350 597020 543922
rect 596400 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597020 526350
rect 596400 526226 597020 526294
rect 596400 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597020 526226
rect 596400 526102 597020 526170
rect 596400 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597020 526102
rect 596400 525978 597020 526046
rect 596400 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597020 525978
rect 596400 508350 597020 525922
rect 596400 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597020 508350
rect 596400 508226 597020 508294
rect 596400 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597020 508226
rect 596400 508102 597020 508170
rect 596400 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597020 508102
rect 596400 507978 597020 508046
rect 596400 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597020 507978
rect 596400 490350 597020 507922
rect 596400 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597020 490350
rect 596400 490226 597020 490294
rect 596400 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597020 490226
rect 596400 490102 597020 490170
rect 596400 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597020 490102
rect 596400 489978 597020 490046
rect 596400 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597020 489978
rect 596400 472350 597020 489922
rect 596400 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597020 472350
rect 596400 472226 597020 472294
rect 596400 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597020 472226
rect 596400 472102 597020 472170
rect 596400 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597020 472102
rect 596400 471978 597020 472046
rect 596400 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597020 471978
rect 596400 454350 597020 471922
rect 596400 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597020 454350
rect 596400 454226 597020 454294
rect 596400 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597020 454226
rect 596400 454102 597020 454170
rect 596400 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597020 454102
rect 596400 453978 597020 454046
rect 596400 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597020 453978
rect 596400 436350 597020 453922
rect 596400 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597020 436350
rect 596400 436226 597020 436294
rect 596400 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597020 436226
rect 596400 436102 597020 436170
rect 596400 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597020 436102
rect 596400 435978 597020 436046
rect 596400 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597020 435978
rect 596400 418350 597020 435922
rect 596400 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597020 418350
rect 596400 418226 597020 418294
rect 596400 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597020 418226
rect 596400 418102 597020 418170
rect 596400 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597020 418102
rect 596400 417978 597020 418046
rect 596400 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597020 417978
rect 596400 400350 597020 417922
rect 596400 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597020 400350
rect 596400 400226 597020 400294
rect 596400 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597020 400226
rect 596400 400102 597020 400170
rect 596400 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597020 400102
rect 596400 399978 597020 400046
rect 596400 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597020 399978
rect 596400 382350 597020 399922
rect 596400 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597020 382350
rect 596400 382226 597020 382294
rect 596400 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597020 382226
rect 596400 382102 597020 382170
rect 596400 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597020 382102
rect 596400 381978 597020 382046
rect 596400 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597020 381978
rect 596400 364350 597020 381922
rect 596400 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597020 364350
rect 596400 364226 597020 364294
rect 596400 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597020 364226
rect 596400 364102 597020 364170
rect 596400 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597020 364102
rect 596400 363978 597020 364046
rect 596400 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597020 363978
rect 596400 346350 597020 363922
rect 596400 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597020 346350
rect 596400 346226 597020 346294
rect 596400 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597020 346226
rect 596400 346102 597020 346170
rect 596400 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597020 346102
rect 596400 345978 597020 346046
rect 596400 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597020 345978
rect 596400 328350 597020 345922
rect 596400 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597020 328350
rect 596400 328226 597020 328294
rect 596400 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597020 328226
rect 596400 328102 597020 328170
rect 596400 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597020 328102
rect 596400 327978 597020 328046
rect 596400 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597020 327978
rect 596400 310350 597020 327922
rect 596400 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597020 310350
rect 596400 310226 597020 310294
rect 596400 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597020 310226
rect 596400 310102 597020 310170
rect 596400 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597020 310102
rect 596400 309978 597020 310046
rect 596400 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597020 309978
rect 596400 292350 597020 309922
rect 596400 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597020 292350
rect 596400 292226 597020 292294
rect 596400 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597020 292226
rect 596400 292102 597020 292170
rect 596400 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597020 292102
rect 596400 291978 597020 292046
rect 596400 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597020 291978
rect 596400 274350 597020 291922
rect 596400 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597020 274350
rect 596400 274226 597020 274294
rect 596400 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597020 274226
rect 596400 274102 597020 274170
rect 596400 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597020 274102
rect 596400 273978 597020 274046
rect 596400 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597020 273978
rect 596400 256350 597020 273922
rect 596400 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597020 256350
rect 596400 256226 597020 256294
rect 596400 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597020 256226
rect 596400 256102 597020 256170
rect 596400 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597020 256102
rect 596400 255978 597020 256046
rect 596400 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597020 255978
rect 596400 238350 597020 255922
rect 596400 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597020 238350
rect 596400 238226 597020 238294
rect 596400 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597020 238226
rect 596400 238102 597020 238170
rect 596400 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597020 238102
rect 596400 237978 597020 238046
rect 596400 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597020 237978
rect 596400 220350 597020 237922
rect 596400 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597020 220350
rect 596400 220226 597020 220294
rect 596400 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597020 220226
rect 596400 220102 597020 220170
rect 596400 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597020 220102
rect 596400 219978 597020 220046
rect 596400 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597020 219978
rect 596400 202350 597020 219922
rect 596400 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597020 202350
rect 596400 202226 597020 202294
rect 596400 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597020 202226
rect 596400 202102 597020 202170
rect 596400 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597020 202102
rect 596400 201978 597020 202046
rect 596400 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597020 201978
rect 596400 184350 597020 201922
rect 596400 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597020 184350
rect 596400 184226 597020 184294
rect 596400 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597020 184226
rect 596400 184102 597020 184170
rect 596400 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597020 184102
rect 596400 183978 597020 184046
rect 596400 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597020 183978
rect 596400 166350 597020 183922
rect 596400 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597020 166350
rect 596400 166226 597020 166294
rect 596400 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597020 166226
rect 596400 166102 597020 166170
rect 596400 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597020 166102
rect 596400 165978 597020 166046
rect 596400 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597020 165978
rect 596400 148350 597020 165922
rect 596400 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597020 148350
rect 596400 148226 597020 148294
rect 596400 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597020 148226
rect 596400 148102 597020 148170
rect 596400 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597020 148102
rect 596400 147978 597020 148046
rect 596400 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597020 147978
rect 596400 130350 597020 147922
rect 596400 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597020 130350
rect 596400 130226 597020 130294
rect 596400 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597020 130226
rect 596400 130102 597020 130170
rect 596400 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597020 130102
rect 596400 129978 597020 130046
rect 596400 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597020 129978
rect 596400 112350 597020 129922
rect 596400 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597020 112350
rect 596400 112226 597020 112294
rect 596400 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597020 112226
rect 596400 112102 597020 112170
rect 596400 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597020 112102
rect 596400 111978 597020 112046
rect 596400 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597020 111978
rect 596400 94350 597020 111922
rect 596400 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597020 94350
rect 596400 94226 597020 94294
rect 596400 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597020 94226
rect 596400 94102 597020 94170
rect 596400 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597020 94102
rect 596400 93978 597020 94046
rect 596400 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597020 93978
rect 596400 76350 597020 93922
rect 596400 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597020 76350
rect 596400 76226 597020 76294
rect 596400 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597020 76226
rect 596400 76102 597020 76170
rect 596400 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597020 76102
rect 596400 75978 597020 76046
rect 596400 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597020 75978
rect 596400 58350 597020 75922
rect 596400 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597020 58350
rect 596400 58226 597020 58294
rect 596400 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597020 58226
rect 596400 58102 597020 58170
rect 596400 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597020 58102
rect 596400 57978 597020 58046
rect 596400 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597020 57978
rect 596400 40350 597020 57922
rect 596400 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597020 40350
rect 596400 40226 597020 40294
rect 596400 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597020 40226
rect 596400 40102 597020 40170
rect 596400 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597020 40102
rect 596400 39978 597020 40046
rect 596400 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597020 39978
rect 596400 22350 597020 39922
rect 596400 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597020 22350
rect 596400 22226 597020 22294
rect 596400 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597020 22226
rect 596400 22102 597020 22170
rect 596400 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597020 22102
rect 596400 21978 597020 22046
rect 596400 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597020 21978
rect 596400 4350 597020 21922
rect 596400 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597020 4350
rect 596400 4226 597020 4294
rect 596400 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597020 4226
rect 596400 4102 597020 4170
rect 596400 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597020 4102
rect 596400 3978 597020 4046
rect 596400 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597020 3978
rect 596400 -160 597020 3922
rect 596400 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect 596400 -284 597020 -216
rect 596400 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect 596400 -408 597020 -340
rect 596400 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect 596400 -532 597020 -464
rect 596400 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect 596400 -684 597020 -588
rect 597360 586350 597980 597744
rect 597360 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect 597360 586226 597980 586294
rect 597360 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect 597360 586102 597980 586170
rect 597360 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect 597360 585978 597980 586046
rect 597360 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect 597360 568350 597980 585922
rect 597360 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect 597360 568226 597980 568294
rect 597360 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect 597360 568102 597980 568170
rect 597360 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect 597360 567978 597980 568046
rect 597360 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect 597360 550350 597980 567922
rect 597360 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect 597360 550226 597980 550294
rect 597360 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect 597360 550102 597980 550170
rect 597360 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect 597360 549978 597980 550046
rect 597360 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect 597360 532350 597980 549922
rect 597360 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect 597360 532226 597980 532294
rect 597360 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect 597360 532102 597980 532170
rect 597360 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect 597360 531978 597980 532046
rect 597360 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect 597360 514350 597980 531922
rect 597360 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect 597360 514226 597980 514294
rect 597360 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect 597360 514102 597980 514170
rect 597360 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect 597360 513978 597980 514046
rect 597360 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect 597360 496350 597980 513922
rect 597360 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect 597360 496226 597980 496294
rect 597360 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect 597360 496102 597980 496170
rect 597360 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect 597360 495978 597980 496046
rect 597360 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect 597360 478350 597980 495922
rect 597360 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect 597360 478226 597980 478294
rect 597360 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect 597360 478102 597980 478170
rect 597360 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect 597360 477978 597980 478046
rect 597360 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect 597360 460350 597980 477922
rect 597360 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect 597360 460226 597980 460294
rect 597360 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect 597360 460102 597980 460170
rect 597360 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect 597360 459978 597980 460046
rect 597360 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect 597360 442350 597980 459922
rect 597360 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect 597360 442226 597980 442294
rect 597360 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect 597360 442102 597980 442170
rect 597360 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect 597360 441978 597980 442046
rect 597360 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect 597360 424350 597980 441922
rect 597360 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect 597360 424226 597980 424294
rect 597360 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect 597360 424102 597980 424170
rect 597360 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect 597360 423978 597980 424046
rect 597360 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect 597360 406350 597980 423922
rect 597360 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect 597360 406226 597980 406294
rect 597360 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect 597360 406102 597980 406170
rect 597360 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect 597360 405978 597980 406046
rect 597360 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect 597360 388350 597980 405922
rect 597360 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect 597360 388226 597980 388294
rect 597360 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect 597360 388102 597980 388170
rect 597360 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect 597360 387978 597980 388046
rect 597360 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect 597360 370350 597980 387922
rect 597360 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect 597360 370226 597980 370294
rect 597360 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect 597360 370102 597980 370170
rect 597360 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect 597360 369978 597980 370046
rect 597360 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect 597360 352350 597980 369922
rect 597360 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect 597360 352226 597980 352294
rect 597360 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect 597360 352102 597980 352170
rect 597360 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect 597360 351978 597980 352046
rect 597360 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect 597360 334350 597980 351922
rect 597360 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect 597360 334226 597980 334294
rect 597360 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect 597360 334102 597980 334170
rect 597360 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect 597360 333978 597980 334046
rect 597360 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect 597360 316350 597980 333922
rect 597360 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect 597360 316226 597980 316294
rect 597360 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect 597360 316102 597980 316170
rect 597360 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect 597360 315978 597980 316046
rect 597360 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect 597360 298350 597980 315922
rect 597360 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect 597360 298226 597980 298294
rect 597360 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect 597360 298102 597980 298170
rect 597360 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect 597360 297978 597980 298046
rect 597360 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect 597360 280350 597980 297922
rect 597360 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect 597360 280226 597980 280294
rect 597360 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect 597360 280102 597980 280170
rect 597360 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect 597360 279978 597980 280046
rect 597360 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect 597360 262350 597980 279922
rect 597360 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect 597360 262226 597980 262294
rect 597360 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect 597360 262102 597980 262170
rect 597360 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect 597360 261978 597980 262046
rect 597360 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect 597360 244350 597980 261922
rect 597360 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect 597360 244226 597980 244294
rect 597360 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect 597360 244102 597980 244170
rect 597360 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect 597360 243978 597980 244046
rect 597360 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect 597360 226350 597980 243922
rect 597360 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect 597360 226226 597980 226294
rect 597360 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect 597360 226102 597980 226170
rect 597360 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect 597360 225978 597980 226046
rect 597360 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect 597360 208350 597980 225922
rect 597360 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect 597360 208226 597980 208294
rect 597360 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect 597360 208102 597980 208170
rect 597360 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect 597360 207978 597980 208046
rect 597360 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect 597360 190350 597980 207922
rect 597360 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect 597360 190226 597980 190294
rect 597360 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect 597360 190102 597980 190170
rect 597360 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect 597360 189978 597980 190046
rect 597360 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect 597360 172350 597980 189922
rect 597360 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect 597360 172226 597980 172294
rect 597360 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect 597360 172102 597980 172170
rect 597360 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect 597360 171978 597980 172046
rect 597360 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect 597360 154350 597980 171922
rect 597360 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect 597360 154226 597980 154294
rect 597360 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect 597360 154102 597980 154170
rect 597360 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect 597360 153978 597980 154046
rect 597360 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect 597360 136350 597980 153922
rect 597360 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect 597360 136226 597980 136294
rect 597360 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect 597360 136102 597980 136170
rect 597360 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect 597360 135978 597980 136046
rect 597360 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect 597360 118350 597980 135922
rect 597360 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect 597360 118226 597980 118294
rect 597360 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect 597360 118102 597980 118170
rect 597360 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect 597360 117978 597980 118046
rect 597360 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect 597360 100350 597980 117922
rect 597360 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect 597360 100226 597980 100294
rect 597360 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect 597360 100102 597980 100170
rect 597360 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect 597360 99978 597980 100046
rect 597360 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect 597360 82350 597980 99922
rect 597360 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect 597360 82226 597980 82294
rect 597360 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect 597360 82102 597980 82170
rect 597360 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect 597360 81978 597980 82046
rect 597360 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect 597360 64350 597980 81922
rect 597360 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect 597360 64226 597980 64294
rect 597360 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect 597360 64102 597980 64170
rect 597360 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect 597360 63978 597980 64046
rect 597360 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect 597360 46350 597980 63922
rect 597360 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect 597360 46226 597980 46294
rect 597360 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect 597360 46102 597980 46170
rect 597360 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect 597360 45978 597980 46046
rect 597360 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect 597360 28350 597980 45922
rect 597360 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect 597360 28226 597980 28294
rect 597360 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect 597360 28102 597980 28170
rect 597360 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect 597360 27978 597980 28046
rect 597360 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect 597360 10350 597980 27922
rect 597360 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect 597360 10226 597980 10294
rect 597360 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect 597360 10102 597980 10170
rect 597360 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect 597360 9978 597980 10046
rect 597360 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect 592818 -1176 592914 -1120
rect 592970 -1176 593038 -1120
rect 593094 -1176 593162 -1120
rect 593218 -1176 593286 -1120
rect 593342 -1176 593438 -1120
rect 592818 -1244 593438 -1176
rect 592818 -1300 592914 -1244
rect 592970 -1300 593038 -1244
rect 593094 -1300 593162 -1244
rect 593218 -1300 593286 -1244
rect 593342 -1300 593438 -1244
rect 592818 -1368 593438 -1300
rect 592818 -1424 592914 -1368
rect 592970 -1424 593038 -1368
rect 593094 -1424 593162 -1368
rect 593218 -1424 593286 -1368
rect 593342 -1424 593438 -1368
rect 592818 -1492 593438 -1424
rect 592818 -1548 592914 -1492
rect 592970 -1548 593038 -1492
rect 593094 -1548 593162 -1492
rect 593218 -1548 593286 -1492
rect 593342 -1548 593438 -1492
rect 592818 -1644 593438 -1548
rect 597360 -1120 597980 9922
rect 597360 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect 597360 -1244 597980 -1176
rect 597360 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect 597360 -1368 597980 -1300
rect 597360 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect 597360 -1492 597980 -1424
rect 597360 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect 597360 -1644 597980 -1548
<< via4 >>
rect -1820 598116 -1764 598172
rect -1696 598116 -1640 598172
rect -1572 598116 -1516 598172
rect -1448 598116 -1392 598172
rect -1820 597992 -1764 598048
rect -1696 597992 -1640 598048
rect -1572 597992 -1516 598048
rect -1448 597992 -1392 598048
rect -1820 597868 -1764 597924
rect -1696 597868 -1640 597924
rect -1572 597868 -1516 597924
rect -1448 597868 -1392 597924
rect -1820 597744 -1764 597800
rect -1696 597744 -1640 597800
rect -1572 597744 -1516 597800
rect -1448 597744 -1392 597800
rect -1820 586294 -1764 586350
rect -1696 586294 -1640 586350
rect -1572 586294 -1516 586350
rect -1448 586294 -1392 586350
rect -1820 586170 -1764 586226
rect -1696 586170 -1640 586226
rect -1572 586170 -1516 586226
rect -1448 586170 -1392 586226
rect -1820 586046 -1764 586102
rect -1696 586046 -1640 586102
rect -1572 586046 -1516 586102
rect -1448 586046 -1392 586102
rect -1820 585922 -1764 585978
rect -1696 585922 -1640 585978
rect -1572 585922 -1516 585978
rect -1448 585922 -1392 585978
rect -1820 568294 -1764 568350
rect -1696 568294 -1640 568350
rect -1572 568294 -1516 568350
rect -1448 568294 -1392 568350
rect -1820 568170 -1764 568226
rect -1696 568170 -1640 568226
rect -1572 568170 -1516 568226
rect -1448 568170 -1392 568226
rect -1820 568046 -1764 568102
rect -1696 568046 -1640 568102
rect -1572 568046 -1516 568102
rect -1448 568046 -1392 568102
rect -1820 567922 -1764 567978
rect -1696 567922 -1640 567978
rect -1572 567922 -1516 567978
rect -1448 567922 -1392 567978
rect -1820 550294 -1764 550350
rect -1696 550294 -1640 550350
rect -1572 550294 -1516 550350
rect -1448 550294 -1392 550350
rect -1820 550170 -1764 550226
rect -1696 550170 -1640 550226
rect -1572 550170 -1516 550226
rect -1448 550170 -1392 550226
rect -1820 550046 -1764 550102
rect -1696 550046 -1640 550102
rect -1572 550046 -1516 550102
rect -1448 550046 -1392 550102
rect -1820 549922 -1764 549978
rect -1696 549922 -1640 549978
rect -1572 549922 -1516 549978
rect -1448 549922 -1392 549978
rect -1820 532294 -1764 532350
rect -1696 532294 -1640 532350
rect -1572 532294 -1516 532350
rect -1448 532294 -1392 532350
rect -1820 532170 -1764 532226
rect -1696 532170 -1640 532226
rect -1572 532170 -1516 532226
rect -1448 532170 -1392 532226
rect -1820 532046 -1764 532102
rect -1696 532046 -1640 532102
rect -1572 532046 -1516 532102
rect -1448 532046 -1392 532102
rect -1820 531922 -1764 531978
rect -1696 531922 -1640 531978
rect -1572 531922 -1516 531978
rect -1448 531922 -1392 531978
rect -1820 514294 -1764 514350
rect -1696 514294 -1640 514350
rect -1572 514294 -1516 514350
rect -1448 514294 -1392 514350
rect -1820 514170 -1764 514226
rect -1696 514170 -1640 514226
rect -1572 514170 -1516 514226
rect -1448 514170 -1392 514226
rect -1820 514046 -1764 514102
rect -1696 514046 -1640 514102
rect -1572 514046 -1516 514102
rect -1448 514046 -1392 514102
rect -1820 513922 -1764 513978
rect -1696 513922 -1640 513978
rect -1572 513922 -1516 513978
rect -1448 513922 -1392 513978
rect -1820 496294 -1764 496350
rect -1696 496294 -1640 496350
rect -1572 496294 -1516 496350
rect -1448 496294 -1392 496350
rect -1820 496170 -1764 496226
rect -1696 496170 -1640 496226
rect -1572 496170 -1516 496226
rect -1448 496170 -1392 496226
rect -1820 496046 -1764 496102
rect -1696 496046 -1640 496102
rect -1572 496046 -1516 496102
rect -1448 496046 -1392 496102
rect -1820 495922 -1764 495978
rect -1696 495922 -1640 495978
rect -1572 495922 -1516 495978
rect -1448 495922 -1392 495978
rect -1820 478294 -1764 478350
rect -1696 478294 -1640 478350
rect -1572 478294 -1516 478350
rect -1448 478294 -1392 478350
rect -1820 478170 -1764 478226
rect -1696 478170 -1640 478226
rect -1572 478170 -1516 478226
rect -1448 478170 -1392 478226
rect -1820 478046 -1764 478102
rect -1696 478046 -1640 478102
rect -1572 478046 -1516 478102
rect -1448 478046 -1392 478102
rect -1820 477922 -1764 477978
rect -1696 477922 -1640 477978
rect -1572 477922 -1516 477978
rect -1448 477922 -1392 477978
rect -1820 460294 -1764 460350
rect -1696 460294 -1640 460350
rect -1572 460294 -1516 460350
rect -1448 460294 -1392 460350
rect -1820 460170 -1764 460226
rect -1696 460170 -1640 460226
rect -1572 460170 -1516 460226
rect -1448 460170 -1392 460226
rect -1820 460046 -1764 460102
rect -1696 460046 -1640 460102
rect -1572 460046 -1516 460102
rect -1448 460046 -1392 460102
rect -1820 459922 -1764 459978
rect -1696 459922 -1640 459978
rect -1572 459922 -1516 459978
rect -1448 459922 -1392 459978
rect -1820 442294 -1764 442350
rect -1696 442294 -1640 442350
rect -1572 442294 -1516 442350
rect -1448 442294 -1392 442350
rect -1820 442170 -1764 442226
rect -1696 442170 -1640 442226
rect -1572 442170 -1516 442226
rect -1448 442170 -1392 442226
rect -1820 442046 -1764 442102
rect -1696 442046 -1640 442102
rect -1572 442046 -1516 442102
rect -1448 442046 -1392 442102
rect -1820 441922 -1764 441978
rect -1696 441922 -1640 441978
rect -1572 441922 -1516 441978
rect -1448 441922 -1392 441978
rect -1820 424294 -1764 424350
rect -1696 424294 -1640 424350
rect -1572 424294 -1516 424350
rect -1448 424294 -1392 424350
rect -1820 424170 -1764 424226
rect -1696 424170 -1640 424226
rect -1572 424170 -1516 424226
rect -1448 424170 -1392 424226
rect -1820 424046 -1764 424102
rect -1696 424046 -1640 424102
rect -1572 424046 -1516 424102
rect -1448 424046 -1392 424102
rect -1820 423922 -1764 423978
rect -1696 423922 -1640 423978
rect -1572 423922 -1516 423978
rect -1448 423922 -1392 423978
rect -1820 406294 -1764 406350
rect -1696 406294 -1640 406350
rect -1572 406294 -1516 406350
rect -1448 406294 -1392 406350
rect -1820 406170 -1764 406226
rect -1696 406170 -1640 406226
rect -1572 406170 -1516 406226
rect -1448 406170 -1392 406226
rect -1820 406046 -1764 406102
rect -1696 406046 -1640 406102
rect -1572 406046 -1516 406102
rect -1448 406046 -1392 406102
rect -1820 405922 -1764 405978
rect -1696 405922 -1640 405978
rect -1572 405922 -1516 405978
rect -1448 405922 -1392 405978
rect -1820 388294 -1764 388350
rect -1696 388294 -1640 388350
rect -1572 388294 -1516 388350
rect -1448 388294 -1392 388350
rect -1820 388170 -1764 388226
rect -1696 388170 -1640 388226
rect -1572 388170 -1516 388226
rect -1448 388170 -1392 388226
rect -1820 388046 -1764 388102
rect -1696 388046 -1640 388102
rect -1572 388046 -1516 388102
rect -1448 388046 -1392 388102
rect -1820 387922 -1764 387978
rect -1696 387922 -1640 387978
rect -1572 387922 -1516 387978
rect -1448 387922 -1392 387978
rect -1820 370294 -1764 370350
rect -1696 370294 -1640 370350
rect -1572 370294 -1516 370350
rect -1448 370294 -1392 370350
rect -1820 370170 -1764 370226
rect -1696 370170 -1640 370226
rect -1572 370170 -1516 370226
rect -1448 370170 -1392 370226
rect -1820 370046 -1764 370102
rect -1696 370046 -1640 370102
rect -1572 370046 -1516 370102
rect -1448 370046 -1392 370102
rect -1820 369922 -1764 369978
rect -1696 369922 -1640 369978
rect -1572 369922 -1516 369978
rect -1448 369922 -1392 369978
rect -1820 352294 -1764 352350
rect -1696 352294 -1640 352350
rect -1572 352294 -1516 352350
rect -1448 352294 -1392 352350
rect -1820 352170 -1764 352226
rect -1696 352170 -1640 352226
rect -1572 352170 -1516 352226
rect -1448 352170 -1392 352226
rect -1820 352046 -1764 352102
rect -1696 352046 -1640 352102
rect -1572 352046 -1516 352102
rect -1448 352046 -1392 352102
rect -1820 351922 -1764 351978
rect -1696 351922 -1640 351978
rect -1572 351922 -1516 351978
rect -1448 351922 -1392 351978
rect -1820 334294 -1764 334350
rect -1696 334294 -1640 334350
rect -1572 334294 -1516 334350
rect -1448 334294 -1392 334350
rect -1820 334170 -1764 334226
rect -1696 334170 -1640 334226
rect -1572 334170 -1516 334226
rect -1448 334170 -1392 334226
rect -1820 334046 -1764 334102
rect -1696 334046 -1640 334102
rect -1572 334046 -1516 334102
rect -1448 334046 -1392 334102
rect -1820 333922 -1764 333978
rect -1696 333922 -1640 333978
rect -1572 333922 -1516 333978
rect -1448 333922 -1392 333978
rect -1820 316294 -1764 316350
rect -1696 316294 -1640 316350
rect -1572 316294 -1516 316350
rect -1448 316294 -1392 316350
rect -1820 316170 -1764 316226
rect -1696 316170 -1640 316226
rect -1572 316170 -1516 316226
rect -1448 316170 -1392 316226
rect -1820 316046 -1764 316102
rect -1696 316046 -1640 316102
rect -1572 316046 -1516 316102
rect -1448 316046 -1392 316102
rect -1820 315922 -1764 315978
rect -1696 315922 -1640 315978
rect -1572 315922 -1516 315978
rect -1448 315922 -1392 315978
rect -1820 298294 -1764 298350
rect -1696 298294 -1640 298350
rect -1572 298294 -1516 298350
rect -1448 298294 -1392 298350
rect -1820 298170 -1764 298226
rect -1696 298170 -1640 298226
rect -1572 298170 -1516 298226
rect -1448 298170 -1392 298226
rect -1820 298046 -1764 298102
rect -1696 298046 -1640 298102
rect -1572 298046 -1516 298102
rect -1448 298046 -1392 298102
rect -1820 297922 -1764 297978
rect -1696 297922 -1640 297978
rect -1572 297922 -1516 297978
rect -1448 297922 -1392 297978
rect -1820 280294 -1764 280350
rect -1696 280294 -1640 280350
rect -1572 280294 -1516 280350
rect -1448 280294 -1392 280350
rect -1820 280170 -1764 280226
rect -1696 280170 -1640 280226
rect -1572 280170 -1516 280226
rect -1448 280170 -1392 280226
rect -1820 280046 -1764 280102
rect -1696 280046 -1640 280102
rect -1572 280046 -1516 280102
rect -1448 280046 -1392 280102
rect -1820 279922 -1764 279978
rect -1696 279922 -1640 279978
rect -1572 279922 -1516 279978
rect -1448 279922 -1392 279978
rect -1820 262294 -1764 262350
rect -1696 262294 -1640 262350
rect -1572 262294 -1516 262350
rect -1448 262294 -1392 262350
rect -1820 262170 -1764 262226
rect -1696 262170 -1640 262226
rect -1572 262170 -1516 262226
rect -1448 262170 -1392 262226
rect -1820 262046 -1764 262102
rect -1696 262046 -1640 262102
rect -1572 262046 -1516 262102
rect -1448 262046 -1392 262102
rect -1820 261922 -1764 261978
rect -1696 261922 -1640 261978
rect -1572 261922 -1516 261978
rect -1448 261922 -1392 261978
rect -1820 244294 -1764 244350
rect -1696 244294 -1640 244350
rect -1572 244294 -1516 244350
rect -1448 244294 -1392 244350
rect -1820 244170 -1764 244226
rect -1696 244170 -1640 244226
rect -1572 244170 -1516 244226
rect -1448 244170 -1392 244226
rect -1820 244046 -1764 244102
rect -1696 244046 -1640 244102
rect -1572 244046 -1516 244102
rect -1448 244046 -1392 244102
rect -1820 243922 -1764 243978
rect -1696 243922 -1640 243978
rect -1572 243922 -1516 243978
rect -1448 243922 -1392 243978
rect -1820 226294 -1764 226350
rect -1696 226294 -1640 226350
rect -1572 226294 -1516 226350
rect -1448 226294 -1392 226350
rect -1820 226170 -1764 226226
rect -1696 226170 -1640 226226
rect -1572 226170 -1516 226226
rect -1448 226170 -1392 226226
rect -1820 226046 -1764 226102
rect -1696 226046 -1640 226102
rect -1572 226046 -1516 226102
rect -1448 226046 -1392 226102
rect -1820 225922 -1764 225978
rect -1696 225922 -1640 225978
rect -1572 225922 -1516 225978
rect -1448 225922 -1392 225978
rect -1820 208294 -1764 208350
rect -1696 208294 -1640 208350
rect -1572 208294 -1516 208350
rect -1448 208294 -1392 208350
rect -1820 208170 -1764 208226
rect -1696 208170 -1640 208226
rect -1572 208170 -1516 208226
rect -1448 208170 -1392 208226
rect -1820 208046 -1764 208102
rect -1696 208046 -1640 208102
rect -1572 208046 -1516 208102
rect -1448 208046 -1392 208102
rect -1820 207922 -1764 207978
rect -1696 207922 -1640 207978
rect -1572 207922 -1516 207978
rect -1448 207922 -1392 207978
rect -1820 190294 -1764 190350
rect -1696 190294 -1640 190350
rect -1572 190294 -1516 190350
rect -1448 190294 -1392 190350
rect -1820 190170 -1764 190226
rect -1696 190170 -1640 190226
rect -1572 190170 -1516 190226
rect -1448 190170 -1392 190226
rect -1820 190046 -1764 190102
rect -1696 190046 -1640 190102
rect -1572 190046 -1516 190102
rect -1448 190046 -1392 190102
rect -1820 189922 -1764 189978
rect -1696 189922 -1640 189978
rect -1572 189922 -1516 189978
rect -1448 189922 -1392 189978
rect -1820 172294 -1764 172350
rect -1696 172294 -1640 172350
rect -1572 172294 -1516 172350
rect -1448 172294 -1392 172350
rect -1820 172170 -1764 172226
rect -1696 172170 -1640 172226
rect -1572 172170 -1516 172226
rect -1448 172170 -1392 172226
rect -1820 172046 -1764 172102
rect -1696 172046 -1640 172102
rect -1572 172046 -1516 172102
rect -1448 172046 -1392 172102
rect -1820 171922 -1764 171978
rect -1696 171922 -1640 171978
rect -1572 171922 -1516 171978
rect -1448 171922 -1392 171978
rect -1820 154294 -1764 154350
rect -1696 154294 -1640 154350
rect -1572 154294 -1516 154350
rect -1448 154294 -1392 154350
rect -1820 154170 -1764 154226
rect -1696 154170 -1640 154226
rect -1572 154170 -1516 154226
rect -1448 154170 -1392 154226
rect -1820 154046 -1764 154102
rect -1696 154046 -1640 154102
rect -1572 154046 -1516 154102
rect -1448 154046 -1392 154102
rect -1820 153922 -1764 153978
rect -1696 153922 -1640 153978
rect -1572 153922 -1516 153978
rect -1448 153922 -1392 153978
rect -1820 136294 -1764 136350
rect -1696 136294 -1640 136350
rect -1572 136294 -1516 136350
rect -1448 136294 -1392 136350
rect -1820 136170 -1764 136226
rect -1696 136170 -1640 136226
rect -1572 136170 -1516 136226
rect -1448 136170 -1392 136226
rect -1820 136046 -1764 136102
rect -1696 136046 -1640 136102
rect -1572 136046 -1516 136102
rect -1448 136046 -1392 136102
rect -1820 135922 -1764 135978
rect -1696 135922 -1640 135978
rect -1572 135922 -1516 135978
rect -1448 135922 -1392 135978
rect -1820 118294 -1764 118350
rect -1696 118294 -1640 118350
rect -1572 118294 -1516 118350
rect -1448 118294 -1392 118350
rect -1820 118170 -1764 118226
rect -1696 118170 -1640 118226
rect -1572 118170 -1516 118226
rect -1448 118170 -1392 118226
rect -1820 118046 -1764 118102
rect -1696 118046 -1640 118102
rect -1572 118046 -1516 118102
rect -1448 118046 -1392 118102
rect -1820 117922 -1764 117978
rect -1696 117922 -1640 117978
rect -1572 117922 -1516 117978
rect -1448 117922 -1392 117978
rect -1820 100294 -1764 100350
rect -1696 100294 -1640 100350
rect -1572 100294 -1516 100350
rect -1448 100294 -1392 100350
rect -1820 100170 -1764 100226
rect -1696 100170 -1640 100226
rect -1572 100170 -1516 100226
rect -1448 100170 -1392 100226
rect -1820 100046 -1764 100102
rect -1696 100046 -1640 100102
rect -1572 100046 -1516 100102
rect -1448 100046 -1392 100102
rect -1820 99922 -1764 99978
rect -1696 99922 -1640 99978
rect -1572 99922 -1516 99978
rect -1448 99922 -1392 99978
rect -1820 82294 -1764 82350
rect -1696 82294 -1640 82350
rect -1572 82294 -1516 82350
rect -1448 82294 -1392 82350
rect -1820 82170 -1764 82226
rect -1696 82170 -1640 82226
rect -1572 82170 -1516 82226
rect -1448 82170 -1392 82226
rect -1820 82046 -1764 82102
rect -1696 82046 -1640 82102
rect -1572 82046 -1516 82102
rect -1448 82046 -1392 82102
rect -1820 81922 -1764 81978
rect -1696 81922 -1640 81978
rect -1572 81922 -1516 81978
rect -1448 81922 -1392 81978
rect -1820 64294 -1764 64350
rect -1696 64294 -1640 64350
rect -1572 64294 -1516 64350
rect -1448 64294 -1392 64350
rect -1820 64170 -1764 64226
rect -1696 64170 -1640 64226
rect -1572 64170 -1516 64226
rect -1448 64170 -1392 64226
rect -1820 64046 -1764 64102
rect -1696 64046 -1640 64102
rect -1572 64046 -1516 64102
rect -1448 64046 -1392 64102
rect -1820 63922 -1764 63978
rect -1696 63922 -1640 63978
rect -1572 63922 -1516 63978
rect -1448 63922 -1392 63978
rect -1820 46294 -1764 46350
rect -1696 46294 -1640 46350
rect -1572 46294 -1516 46350
rect -1448 46294 -1392 46350
rect -1820 46170 -1764 46226
rect -1696 46170 -1640 46226
rect -1572 46170 -1516 46226
rect -1448 46170 -1392 46226
rect -1820 46046 -1764 46102
rect -1696 46046 -1640 46102
rect -1572 46046 -1516 46102
rect -1448 46046 -1392 46102
rect -1820 45922 -1764 45978
rect -1696 45922 -1640 45978
rect -1572 45922 -1516 45978
rect -1448 45922 -1392 45978
rect -1820 28294 -1764 28350
rect -1696 28294 -1640 28350
rect -1572 28294 -1516 28350
rect -1448 28294 -1392 28350
rect -1820 28170 -1764 28226
rect -1696 28170 -1640 28226
rect -1572 28170 -1516 28226
rect -1448 28170 -1392 28226
rect -1820 28046 -1764 28102
rect -1696 28046 -1640 28102
rect -1572 28046 -1516 28102
rect -1448 28046 -1392 28102
rect -1820 27922 -1764 27978
rect -1696 27922 -1640 27978
rect -1572 27922 -1516 27978
rect -1448 27922 -1392 27978
rect -1820 10294 -1764 10350
rect -1696 10294 -1640 10350
rect -1572 10294 -1516 10350
rect -1448 10294 -1392 10350
rect -1820 10170 -1764 10226
rect -1696 10170 -1640 10226
rect -1572 10170 -1516 10226
rect -1448 10170 -1392 10226
rect -1820 10046 -1764 10102
rect -1696 10046 -1640 10102
rect -1572 10046 -1516 10102
rect -1448 10046 -1392 10102
rect -1820 9922 -1764 9978
rect -1696 9922 -1640 9978
rect -1572 9922 -1516 9978
rect -1448 9922 -1392 9978
rect -860 597156 -804 597212
rect -736 597156 -680 597212
rect -612 597156 -556 597212
rect -488 597156 -432 597212
rect -860 597032 -804 597088
rect -736 597032 -680 597088
rect -612 597032 -556 597088
rect -488 597032 -432 597088
rect -860 596908 -804 596964
rect -736 596908 -680 596964
rect -612 596908 -556 596964
rect -488 596908 -432 596964
rect -860 596784 -804 596840
rect -736 596784 -680 596840
rect -612 596784 -556 596840
rect -488 596784 -432 596840
rect 5514 597156 5570 597212
rect 5638 597156 5694 597212
rect 5762 597156 5818 597212
rect 5886 597156 5942 597212
rect 5514 597032 5570 597088
rect 5638 597032 5694 597088
rect 5762 597032 5818 597088
rect 5886 597032 5942 597088
rect 5514 596908 5570 596964
rect 5638 596908 5694 596964
rect 5762 596908 5818 596964
rect 5886 596908 5942 596964
rect 5514 596784 5570 596840
rect 5638 596784 5694 596840
rect 5762 596784 5818 596840
rect 5886 596784 5942 596840
rect -860 580294 -804 580350
rect -736 580294 -680 580350
rect -612 580294 -556 580350
rect -488 580294 -432 580350
rect -860 580170 -804 580226
rect -736 580170 -680 580226
rect -612 580170 -556 580226
rect -488 580170 -432 580226
rect -860 580046 -804 580102
rect -736 580046 -680 580102
rect -612 580046 -556 580102
rect -488 580046 -432 580102
rect -860 579922 -804 579978
rect -736 579922 -680 579978
rect -612 579922 -556 579978
rect -488 579922 -432 579978
rect 9234 598116 9290 598172
rect 9358 598116 9414 598172
rect 9482 598116 9538 598172
rect 9606 598116 9662 598172
rect 9234 597992 9290 598048
rect 9358 597992 9414 598048
rect 9482 597992 9538 598048
rect 9606 597992 9662 598048
rect 9234 597868 9290 597924
rect 9358 597868 9414 597924
rect 9482 597868 9538 597924
rect 9606 597868 9662 597924
rect 9234 597744 9290 597800
rect 9358 597744 9414 597800
rect 9482 597744 9538 597800
rect 9606 597744 9662 597800
rect 9234 586294 9290 586350
rect 9358 586294 9414 586350
rect 9482 586294 9538 586350
rect 9606 586294 9662 586350
rect 9234 586170 9290 586226
rect 9358 586170 9414 586226
rect 9482 586170 9538 586226
rect 9606 586170 9662 586226
rect 9234 586046 9290 586102
rect 9358 586046 9414 586102
rect 9482 586046 9538 586102
rect 9606 586046 9662 586102
rect 9234 585922 9290 585978
rect 9358 585922 9414 585978
rect 9482 585922 9538 585978
rect 9606 585922 9662 585978
rect 39954 598116 40010 598172
rect 40078 598116 40134 598172
rect 40202 598116 40258 598172
rect 40326 598116 40382 598172
rect 39954 597992 40010 598048
rect 40078 597992 40134 598048
rect 40202 597992 40258 598048
rect 40326 597992 40382 598048
rect 39954 597868 40010 597924
rect 40078 597868 40134 597924
rect 40202 597868 40258 597924
rect 40326 597868 40382 597924
rect 39954 597744 40010 597800
rect 40078 597744 40134 597800
rect 40202 597744 40258 597800
rect 40326 597744 40382 597800
rect 39954 586294 40010 586350
rect 40078 586294 40134 586350
rect 40202 586294 40258 586350
rect 40326 586294 40382 586350
rect 39954 586170 40010 586226
rect 40078 586170 40134 586226
rect 40202 586170 40258 586226
rect 40326 586170 40382 586226
rect 39954 586046 40010 586102
rect 40078 586046 40134 586102
rect 40202 586046 40258 586102
rect 40326 586046 40382 586102
rect 39954 585922 40010 585978
rect 40078 585922 40134 585978
rect 40202 585922 40258 585978
rect 40326 585922 40382 585978
rect 70674 598116 70730 598172
rect 70798 598116 70854 598172
rect 70922 598116 70978 598172
rect 71046 598116 71102 598172
rect 70674 597992 70730 598048
rect 70798 597992 70854 598048
rect 70922 597992 70978 598048
rect 71046 597992 71102 598048
rect 70674 597868 70730 597924
rect 70798 597868 70854 597924
rect 70922 597868 70978 597924
rect 71046 597868 71102 597924
rect 70674 597744 70730 597800
rect 70798 597744 70854 597800
rect 70922 597744 70978 597800
rect 71046 597744 71102 597800
rect 70674 586294 70730 586350
rect 70798 586294 70854 586350
rect 70922 586294 70978 586350
rect 71046 586294 71102 586350
rect 70674 586170 70730 586226
rect 70798 586170 70854 586226
rect 70922 586170 70978 586226
rect 71046 586170 71102 586226
rect 70674 586046 70730 586102
rect 70798 586046 70854 586102
rect 70922 586046 70978 586102
rect 71046 586046 71102 586102
rect 70674 585922 70730 585978
rect 70798 585922 70854 585978
rect 70922 585922 70978 585978
rect 71046 585922 71102 585978
rect 101394 598116 101450 598172
rect 101518 598116 101574 598172
rect 101642 598116 101698 598172
rect 101766 598116 101822 598172
rect 101394 597992 101450 598048
rect 101518 597992 101574 598048
rect 101642 597992 101698 598048
rect 101766 597992 101822 598048
rect 101394 597868 101450 597924
rect 101518 597868 101574 597924
rect 101642 597868 101698 597924
rect 101766 597868 101822 597924
rect 101394 597744 101450 597800
rect 101518 597744 101574 597800
rect 101642 597744 101698 597800
rect 101766 597744 101822 597800
rect 101394 586294 101450 586350
rect 101518 586294 101574 586350
rect 101642 586294 101698 586350
rect 101766 586294 101822 586350
rect 101394 586170 101450 586226
rect 101518 586170 101574 586226
rect 101642 586170 101698 586226
rect 101766 586170 101822 586226
rect 101394 586046 101450 586102
rect 101518 586046 101574 586102
rect 101642 586046 101698 586102
rect 101766 586046 101822 586102
rect 101394 585922 101450 585978
rect 101518 585922 101574 585978
rect 101642 585922 101698 585978
rect 101766 585922 101822 585978
rect 132114 598116 132170 598172
rect 132238 598116 132294 598172
rect 132362 598116 132418 598172
rect 132486 598116 132542 598172
rect 132114 597992 132170 598048
rect 132238 597992 132294 598048
rect 132362 597992 132418 598048
rect 132486 597992 132542 598048
rect 132114 597868 132170 597924
rect 132238 597868 132294 597924
rect 132362 597868 132418 597924
rect 132486 597868 132542 597924
rect 132114 597744 132170 597800
rect 132238 597744 132294 597800
rect 132362 597744 132418 597800
rect 132486 597744 132542 597800
rect 132114 586294 132170 586350
rect 132238 586294 132294 586350
rect 132362 586294 132418 586350
rect 132486 586294 132542 586350
rect 132114 586170 132170 586226
rect 132238 586170 132294 586226
rect 132362 586170 132418 586226
rect 132486 586170 132542 586226
rect 132114 586046 132170 586102
rect 132238 586046 132294 586102
rect 132362 586046 132418 586102
rect 132486 586046 132542 586102
rect 132114 585922 132170 585978
rect 132238 585922 132294 585978
rect 132362 585922 132418 585978
rect 132486 585922 132542 585978
rect 162834 598116 162890 598172
rect 162958 598116 163014 598172
rect 163082 598116 163138 598172
rect 163206 598116 163262 598172
rect 162834 597992 162890 598048
rect 162958 597992 163014 598048
rect 163082 597992 163138 598048
rect 163206 597992 163262 598048
rect 162834 597868 162890 597924
rect 162958 597868 163014 597924
rect 163082 597868 163138 597924
rect 163206 597868 163262 597924
rect 162834 597744 162890 597800
rect 162958 597744 163014 597800
rect 163082 597744 163138 597800
rect 163206 597744 163262 597800
rect 162834 586294 162890 586350
rect 162958 586294 163014 586350
rect 163082 586294 163138 586350
rect 163206 586294 163262 586350
rect 162834 586170 162890 586226
rect 162958 586170 163014 586226
rect 163082 586170 163138 586226
rect 163206 586170 163262 586226
rect 162834 586046 162890 586102
rect 162958 586046 163014 586102
rect 163082 586046 163138 586102
rect 163206 586046 163262 586102
rect 162834 585922 162890 585978
rect 162958 585922 163014 585978
rect 163082 585922 163138 585978
rect 163206 585922 163262 585978
rect 193554 598116 193610 598172
rect 193678 598116 193734 598172
rect 193802 598116 193858 598172
rect 193926 598116 193982 598172
rect 193554 597992 193610 598048
rect 193678 597992 193734 598048
rect 193802 597992 193858 598048
rect 193926 597992 193982 598048
rect 193554 597868 193610 597924
rect 193678 597868 193734 597924
rect 193802 597868 193858 597924
rect 193926 597868 193982 597924
rect 193554 597744 193610 597800
rect 193678 597744 193734 597800
rect 193802 597744 193858 597800
rect 193926 597744 193982 597800
rect 193554 586294 193610 586350
rect 193678 586294 193734 586350
rect 193802 586294 193858 586350
rect 193926 586294 193982 586350
rect 193554 586170 193610 586226
rect 193678 586170 193734 586226
rect 193802 586170 193858 586226
rect 193926 586170 193982 586226
rect 193554 586046 193610 586102
rect 193678 586046 193734 586102
rect 193802 586046 193858 586102
rect 193926 586046 193982 586102
rect 193554 585922 193610 585978
rect 193678 585922 193734 585978
rect 193802 585922 193858 585978
rect 193926 585922 193982 585978
rect 224274 598116 224330 598172
rect 224398 598116 224454 598172
rect 224522 598116 224578 598172
rect 224646 598116 224702 598172
rect 224274 597992 224330 598048
rect 224398 597992 224454 598048
rect 224522 597992 224578 598048
rect 224646 597992 224702 598048
rect 224274 597868 224330 597924
rect 224398 597868 224454 597924
rect 224522 597868 224578 597924
rect 224646 597868 224702 597924
rect 224274 597744 224330 597800
rect 224398 597744 224454 597800
rect 224522 597744 224578 597800
rect 224646 597744 224702 597800
rect 224274 586294 224330 586350
rect 224398 586294 224454 586350
rect 224522 586294 224578 586350
rect 224646 586294 224702 586350
rect 224274 586170 224330 586226
rect 224398 586170 224454 586226
rect 224522 586170 224578 586226
rect 224646 586170 224702 586226
rect 224274 586046 224330 586102
rect 224398 586046 224454 586102
rect 224522 586046 224578 586102
rect 224646 586046 224702 586102
rect 224274 585922 224330 585978
rect 224398 585922 224454 585978
rect 224522 585922 224578 585978
rect 224646 585922 224702 585978
rect 254994 598116 255050 598172
rect 255118 598116 255174 598172
rect 255242 598116 255298 598172
rect 255366 598116 255422 598172
rect 254994 597992 255050 598048
rect 255118 597992 255174 598048
rect 255242 597992 255298 598048
rect 255366 597992 255422 598048
rect 254994 597868 255050 597924
rect 255118 597868 255174 597924
rect 255242 597868 255298 597924
rect 255366 597868 255422 597924
rect 254994 597744 255050 597800
rect 255118 597744 255174 597800
rect 255242 597744 255298 597800
rect 255366 597744 255422 597800
rect 254994 586294 255050 586350
rect 255118 586294 255174 586350
rect 255242 586294 255298 586350
rect 255366 586294 255422 586350
rect 254994 586170 255050 586226
rect 255118 586170 255174 586226
rect 255242 586170 255298 586226
rect 255366 586170 255422 586226
rect 254994 586046 255050 586102
rect 255118 586046 255174 586102
rect 255242 586046 255298 586102
rect 255366 586046 255422 586102
rect 254994 585922 255050 585978
rect 255118 585922 255174 585978
rect 255242 585922 255298 585978
rect 255366 585922 255422 585978
rect 285714 598116 285770 598172
rect 285838 598116 285894 598172
rect 285962 598116 286018 598172
rect 286086 598116 286142 598172
rect 285714 597992 285770 598048
rect 285838 597992 285894 598048
rect 285962 597992 286018 598048
rect 286086 597992 286142 598048
rect 285714 597868 285770 597924
rect 285838 597868 285894 597924
rect 285962 597868 286018 597924
rect 286086 597868 286142 597924
rect 285714 597744 285770 597800
rect 285838 597744 285894 597800
rect 285962 597744 286018 597800
rect 286086 597744 286142 597800
rect 285714 586294 285770 586350
rect 285838 586294 285894 586350
rect 285962 586294 286018 586350
rect 286086 586294 286142 586350
rect 285714 586170 285770 586226
rect 285838 586170 285894 586226
rect 285962 586170 286018 586226
rect 286086 586170 286142 586226
rect 285714 586046 285770 586102
rect 285838 586046 285894 586102
rect 285962 586046 286018 586102
rect 286086 586046 286142 586102
rect 285714 585922 285770 585978
rect 285838 585922 285894 585978
rect 285962 585922 286018 585978
rect 286086 585922 286142 585978
rect 316434 598116 316490 598172
rect 316558 598116 316614 598172
rect 316682 598116 316738 598172
rect 316806 598116 316862 598172
rect 316434 597992 316490 598048
rect 316558 597992 316614 598048
rect 316682 597992 316738 598048
rect 316806 597992 316862 598048
rect 316434 597868 316490 597924
rect 316558 597868 316614 597924
rect 316682 597868 316738 597924
rect 316806 597868 316862 597924
rect 316434 597744 316490 597800
rect 316558 597744 316614 597800
rect 316682 597744 316738 597800
rect 316806 597744 316862 597800
rect 316434 586294 316490 586350
rect 316558 586294 316614 586350
rect 316682 586294 316738 586350
rect 316806 586294 316862 586350
rect 316434 586170 316490 586226
rect 316558 586170 316614 586226
rect 316682 586170 316738 586226
rect 316806 586170 316862 586226
rect 316434 586046 316490 586102
rect 316558 586046 316614 586102
rect 316682 586046 316738 586102
rect 316806 586046 316862 586102
rect 316434 585922 316490 585978
rect 316558 585922 316614 585978
rect 316682 585922 316738 585978
rect 316806 585922 316862 585978
rect 347154 598116 347210 598172
rect 347278 598116 347334 598172
rect 347402 598116 347458 598172
rect 347526 598116 347582 598172
rect 347154 597992 347210 598048
rect 347278 597992 347334 598048
rect 347402 597992 347458 598048
rect 347526 597992 347582 598048
rect 347154 597868 347210 597924
rect 347278 597868 347334 597924
rect 347402 597868 347458 597924
rect 347526 597868 347582 597924
rect 347154 597744 347210 597800
rect 347278 597744 347334 597800
rect 347402 597744 347458 597800
rect 347526 597744 347582 597800
rect 347154 586294 347210 586350
rect 347278 586294 347334 586350
rect 347402 586294 347458 586350
rect 347526 586294 347582 586350
rect 347154 586170 347210 586226
rect 347278 586170 347334 586226
rect 347402 586170 347458 586226
rect 347526 586170 347582 586226
rect 347154 586046 347210 586102
rect 347278 586046 347334 586102
rect 347402 586046 347458 586102
rect 347526 586046 347582 586102
rect 347154 585922 347210 585978
rect 347278 585922 347334 585978
rect 347402 585922 347458 585978
rect 347526 585922 347582 585978
rect 377874 598116 377930 598172
rect 377998 598116 378054 598172
rect 378122 598116 378178 598172
rect 378246 598116 378302 598172
rect 377874 597992 377930 598048
rect 377998 597992 378054 598048
rect 378122 597992 378178 598048
rect 378246 597992 378302 598048
rect 377874 597868 377930 597924
rect 377998 597868 378054 597924
rect 378122 597868 378178 597924
rect 378246 597868 378302 597924
rect 377874 597744 377930 597800
rect 377998 597744 378054 597800
rect 378122 597744 378178 597800
rect 378246 597744 378302 597800
rect 377874 586294 377930 586350
rect 377998 586294 378054 586350
rect 378122 586294 378178 586350
rect 378246 586294 378302 586350
rect 377874 586170 377930 586226
rect 377998 586170 378054 586226
rect 378122 586170 378178 586226
rect 378246 586170 378302 586226
rect 377874 586046 377930 586102
rect 377998 586046 378054 586102
rect 378122 586046 378178 586102
rect 378246 586046 378302 586102
rect 377874 585922 377930 585978
rect 377998 585922 378054 585978
rect 378122 585922 378178 585978
rect 378246 585922 378302 585978
rect 408594 598116 408650 598172
rect 408718 598116 408774 598172
rect 408842 598116 408898 598172
rect 408966 598116 409022 598172
rect 408594 597992 408650 598048
rect 408718 597992 408774 598048
rect 408842 597992 408898 598048
rect 408966 597992 409022 598048
rect 408594 597868 408650 597924
rect 408718 597868 408774 597924
rect 408842 597868 408898 597924
rect 408966 597868 409022 597924
rect 408594 597744 408650 597800
rect 408718 597744 408774 597800
rect 408842 597744 408898 597800
rect 408966 597744 409022 597800
rect 408594 586294 408650 586350
rect 408718 586294 408774 586350
rect 408842 586294 408898 586350
rect 408966 586294 409022 586350
rect 408594 586170 408650 586226
rect 408718 586170 408774 586226
rect 408842 586170 408898 586226
rect 408966 586170 409022 586226
rect 408594 586046 408650 586102
rect 408718 586046 408774 586102
rect 408842 586046 408898 586102
rect 408966 586046 409022 586102
rect 408594 585922 408650 585978
rect 408718 585922 408774 585978
rect 408842 585922 408898 585978
rect 408966 585922 409022 585978
rect 439314 598116 439370 598172
rect 439438 598116 439494 598172
rect 439562 598116 439618 598172
rect 439686 598116 439742 598172
rect 439314 597992 439370 598048
rect 439438 597992 439494 598048
rect 439562 597992 439618 598048
rect 439686 597992 439742 598048
rect 439314 597868 439370 597924
rect 439438 597868 439494 597924
rect 439562 597868 439618 597924
rect 439686 597868 439742 597924
rect 439314 597744 439370 597800
rect 439438 597744 439494 597800
rect 439562 597744 439618 597800
rect 439686 597744 439742 597800
rect 439314 586294 439370 586350
rect 439438 586294 439494 586350
rect 439562 586294 439618 586350
rect 439686 586294 439742 586350
rect 439314 586170 439370 586226
rect 439438 586170 439494 586226
rect 439562 586170 439618 586226
rect 439686 586170 439742 586226
rect 439314 586046 439370 586102
rect 439438 586046 439494 586102
rect 439562 586046 439618 586102
rect 439686 586046 439742 586102
rect 439314 585922 439370 585978
rect 439438 585922 439494 585978
rect 439562 585922 439618 585978
rect 439686 585922 439742 585978
rect 470034 598116 470090 598172
rect 470158 598116 470214 598172
rect 470282 598116 470338 598172
rect 470406 598116 470462 598172
rect 470034 597992 470090 598048
rect 470158 597992 470214 598048
rect 470282 597992 470338 598048
rect 470406 597992 470462 598048
rect 470034 597868 470090 597924
rect 470158 597868 470214 597924
rect 470282 597868 470338 597924
rect 470406 597868 470462 597924
rect 470034 597744 470090 597800
rect 470158 597744 470214 597800
rect 470282 597744 470338 597800
rect 470406 597744 470462 597800
rect 470034 586294 470090 586350
rect 470158 586294 470214 586350
rect 470282 586294 470338 586350
rect 470406 586294 470462 586350
rect 470034 586170 470090 586226
rect 470158 586170 470214 586226
rect 470282 586170 470338 586226
rect 470406 586170 470462 586226
rect 470034 586046 470090 586102
rect 470158 586046 470214 586102
rect 470282 586046 470338 586102
rect 470406 586046 470462 586102
rect 470034 585922 470090 585978
rect 470158 585922 470214 585978
rect 470282 585922 470338 585978
rect 470406 585922 470462 585978
rect 500754 598116 500810 598172
rect 500878 598116 500934 598172
rect 501002 598116 501058 598172
rect 501126 598116 501182 598172
rect 500754 597992 500810 598048
rect 500878 597992 500934 598048
rect 501002 597992 501058 598048
rect 501126 597992 501182 598048
rect 500754 597868 500810 597924
rect 500878 597868 500934 597924
rect 501002 597868 501058 597924
rect 501126 597868 501182 597924
rect 500754 597744 500810 597800
rect 500878 597744 500934 597800
rect 501002 597744 501058 597800
rect 501126 597744 501182 597800
rect 500754 586294 500810 586350
rect 500878 586294 500934 586350
rect 501002 586294 501058 586350
rect 501126 586294 501182 586350
rect 500754 586170 500810 586226
rect 500878 586170 500934 586226
rect 501002 586170 501058 586226
rect 501126 586170 501182 586226
rect 500754 586046 500810 586102
rect 500878 586046 500934 586102
rect 501002 586046 501058 586102
rect 501126 586046 501182 586102
rect 500754 585922 500810 585978
rect 500878 585922 500934 585978
rect 501002 585922 501058 585978
rect 501126 585922 501182 585978
rect 531474 598116 531530 598172
rect 531598 598116 531654 598172
rect 531722 598116 531778 598172
rect 531846 598116 531902 598172
rect 531474 597992 531530 598048
rect 531598 597992 531654 598048
rect 531722 597992 531778 598048
rect 531846 597992 531902 598048
rect 531474 597868 531530 597924
rect 531598 597868 531654 597924
rect 531722 597868 531778 597924
rect 531846 597868 531902 597924
rect 531474 597744 531530 597800
rect 531598 597744 531654 597800
rect 531722 597744 531778 597800
rect 531846 597744 531902 597800
rect 531474 586294 531530 586350
rect 531598 586294 531654 586350
rect 531722 586294 531778 586350
rect 531846 586294 531902 586350
rect 531474 586170 531530 586226
rect 531598 586170 531654 586226
rect 531722 586170 531778 586226
rect 531846 586170 531902 586226
rect 531474 586046 531530 586102
rect 531598 586046 531654 586102
rect 531722 586046 531778 586102
rect 531846 586046 531902 586102
rect 531474 585922 531530 585978
rect 531598 585922 531654 585978
rect 531722 585922 531778 585978
rect 531846 585922 531902 585978
rect 562194 598116 562250 598172
rect 562318 598116 562374 598172
rect 562442 598116 562498 598172
rect 562566 598116 562622 598172
rect 562194 597992 562250 598048
rect 562318 597992 562374 598048
rect 562442 597992 562498 598048
rect 562566 597992 562622 598048
rect 562194 597868 562250 597924
rect 562318 597868 562374 597924
rect 562442 597868 562498 597924
rect 562566 597868 562622 597924
rect 562194 597744 562250 597800
rect 562318 597744 562374 597800
rect 562442 597744 562498 597800
rect 562566 597744 562622 597800
rect 562194 586294 562250 586350
rect 562318 586294 562374 586350
rect 562442 586294 562498 586350
rect 562566 586294 562622 586350
rect 562194 586170 562250 586226
rect 562318 586170 562374 586226
rect 562442 586170 562498 586226
rect 562566 586170 562622 586226
rect 562194 586046 562250 586102
rect 562318 586046 562374 586102
rect 562442 586046 562498 586102
rect 562566 586046 562622 586102
rect 562194 585922 562250 585978
rect 562318 585922 562374 585978
rect 562442 585922 562498 585978
rect 562566 585922 562622 585978
rect 589194 597156 589250 597212
rect 589318 597156 589374 597212
rect 589442 597156 589498 597212
rect 589566 597156 589622 597212
rect 589194 597032 589250 597088
rect 589318 597032 589374 597088
rect 589442 597032 589498 597088
rect 589566 597032 589622 597088
rect 589194 596908 589250 596964
rect 589318 596908 589374 596964
rect 589442 596908 589498 596964
rect 589566 596908 589622 596964
rect 589194 596784 589250 596840
rect 589318 596784 589374 596840
rect 589442 596784 589498 596840
rect 589566 596784 589622 596840
rect 5514 580294 5570 580350
rect 5638 580294 5694 580350
rect 5762 580294 5818 580350
rect 5886 580294 5942 580350
rect 5514 580170 5570 580226
rect 5638 580170 5694 580226
rect 5762 580170 5818 580226
rect 5886 580170 5942 580226
rect 5514 580046 5570 580102
rect 5638 580046 5694 580102
rect 5762 580046 5818 580102
rect 5886 580046 5942 580102
rect 5514 579922 5570 579978
rect 5638 579922 5694 579978
rect 5762 579922 5818 579978
rect 5886 579922 5942 579978
rect -860 562294 -804 562350
rect -736 562294 -680 562350
rect -612 562294 -556 562350
rect -488 562294 -432 562350
rect -860 562170 -804 562226
rect -736 562170 -680 562226
rect -612 562170 -556 562226
rect -488 562170 -432 562226
rect -860 562046 -804 562102
rect -736 562046 -680 562102
rect -612 562046 -556 562102
rect -488 562046 -432 562102
rect -860 561922 -804 561978
rect -736 561922 -680 561978
rect -612 561922 -556 561978
rect -488 561922 -432 561978
rect 12518 580294 12574 580350
rect 12642 580294 12698 580350
rect 12518 580170 12574 580226
rect 12642 580170 12698 580226
rect 12518 580046 12574 580102
rect 12642 580046 12698 580102
rect 12518 579922 12574 579978
rect 12642 579922 12698 579978
rect 43238 580294 43294 580350
rect 43362 580294 43418 580350
rect 43238 580170 43294 580226
rect 43362 580170 43418 580226
rect 43238 580046 43294 580102
rect 43362 580046 43418 580102
rect 43238 579922 43294 579978
rect 43362 579922 43418 579978
rect 73958 580294 74014 580350
rect 74082 580294 74138 580350
rect 73958 580170 74014 580226
rect 74082 580170 74138 580226
rect 73958 580046 74014 580102
rect 74082 580046 74138 580102
rect 73958 579922 74014 579978
rect 74082 579922 74138 579978
rect 104678 580294 104734 580350
rect 104802 580294 104858 580350
rect 104678 580170 104734 580226
rect 104802 580170 104858 580226
rect 104678 580046 104734 580102
rect 104802 580046 104858 580102
rect 104678 579922 104734 579978
rect 104802 579922 104858 579978
rect 135398 580294 135454 580350
rect 135522 580294 135578 580350
rect 135398 580170 135454 580226
rect 135522 580170 135578 580226
rect 135398 580046 135454 580102
rect 135522 580046 135578 580102
rect 135398 579922 135454 579978
rect 135522 579922 135578 579978
rect 166118 580294 166174 580350
rect 166242 580294 166298 580350
rect 166118 580170 166174 580226
rect 166242 580170 166298 580226
rect 166118 580046 166174 580102
rect 166242 580046 166298 580102
rect 166118 579922 166174 579978
rect 166242 579922 166298 579978
rect 196838 580294 196894 580350
rect 196962 580294 197018 580350
rect 196838 580170 196894 580226
rect 196962 580170 197018 580226
rect 196838 580046 196894 580102
rect 196962 580046 197018 580102
rect 196838 579922 196894 579978
rect 196962 579922 197018 579978
rect 227558 580294 227614 580350
rect 227682 580294 227738 580350
rect 227558 580170 227614 580226
rect 227682 580170 227738 580226
rect 227558 580046 227614 580102
rect 227682 580046 227738 580102
rect 227558 579922 227614 579978
rect 227682 579922 227738 579978
rect 258278 580294 258334 580350
rect 258402 580294 258458 580350
rect 258278 580170 258334 580226
rect 258402 580170 258458 580226
rect 258278 580046 258334 580102
rect 258402 580046 258458 580102
rect 258278 579922 258334 579978
rect 258402 579922 258458 579978
rect 288998 580294 289054 580350
rect 289122 580294 289178 580350
rect 288998 580170 289054 580226
rect 289122 580170 289178 580226
rect 288998 580046 289054 580102
rect 289122 580046 289178 580102
rect 288998 579922 289054 579978
rect 289122 579922 289178 579978
rect 319718 580294 319774 580350
rect 319842 580294 319898 580350
rect 319718 580170 319774 580226
rect 319842 580170 319898 580226
rect 319718 580046 319774 580102
rect 319842 580046 319898 580102
rect 319718 579922 319774 579978
rect 319842 579922 319898 579978
rect 350438 580294 350494 580350
rect 350562 580294 350618 580350
rect 350438 580170 350494 580226
rect 350562 580170 350618 580226
rect 350438 580046 350494 580102
rect 350562 580046 350618 580102
rect 350438 579922 350494 579978
rect 350562 579922 350618 579978
rect 381158 580294 381214 580350
rect 381282 580294 381338 580350
rect 381158 580170 381214 580226
rect 381282 580170 381338 580226
rect 381158 580046 381214 580102
rect 381282 580046 381338 580102
rect 381158 579922 381214 579978
rect 381282 579922 381338 579978
rect 411878 580294 411934 580350
rect 412002 580294 412058 580350
rect 411878 580170 411934 580226
rect 412002 580170 412058 580226
rect 411878 580046 411934 580102
rect 412002 580046 412058 580102
rect 411878 579922 411934 579978
rect 412002 579922 412058 579978
rect 442598 580294 442654 580350
rect 442722 580294 442778 580350
rect 442598 580170 442654 580226
rect 442722 580170 442778 580226
rect 442598 580046 442654 580102
rect 442722 580046 442778 580102
rect 442598 579922 442654 579978
rect 442722 579922 442778 579978
rect 473318 580294 473374 580350
rect 473442 580294 473498 580350
rect 473318 580170 473374 580226
rect 473442 580170 473498 580226
rect 473318 580046 473374 580102
rect 473442 580046 473498 580102
rect 473318 579922 473374 579978
rect 473442 579922 473498 579978
rect 504038 580294 504094 580350
rect 504162 580294 504218 580350
rect 504038 580170 504094 580226
rect 504162 580170 504218 580226
rect 504038 580046 504094 580102
rect 504162 580046 504218 580102
rect 504038 579922 504094 579978
rect 504162 579922 504218 579978
rect 534758 580294 534814 580350
rect 534882 580294 534938 580350
rect 534758 580170 534814 580226
rect 534882 580170 534938 580226
rect 534758 580046 534814 580102
rect 534882 580046 534938 580102
rect 534758 579922 534814 579978
rect 534882 579922 534938 579978
rect 565478 580294 565534 580350
rect 565602 580294 565658 580350
rect 565478 580170 565534 580226
rect 565602 580170 565658 580226
rect 565478 580046 565534 580102
rect 565602 580046 565658 580102
rect 565478 579922 565534 579978
rect 565602 579922 565658 579978
rect 592914 598116 592970 598172
rect 593038 598116 593094 598172
rect 593162 598116 593218 598172
rect 593286 598116 593342 598172
rect 592914 597992 592970 598048
rect 593038 597992 593094 598048
rect 593162 597992 593218 598048
rect 593286 597992 593342 598048
rect 592914 597868 592970 597924
rect 593038 597868 593094 597924
rect 593162 597868 593218 597924
rect 593286 597868 593342 597924
rect 592914 597744 592970 597800
rect 593038 597744 593094 597800
rect 593162 597744 593218 597800
rect 593286 597744 593342 597800
rect 589194 580294 589250 580350
rect 589318 580294 589374 580350
rect 589442 580294 589498 580350
rect 589566 580294 589622 580350
rect 589194 580170 589250 580226
rect 589318 580170 589374 580226
rect 589442 580170 589498 580226
rect 589566 580170 589622 580226
rect 589194 580046 589250 580102
rect 589318 580046 589374 580102
rect 589442 580046 589498 580102
rect 589566 580046 589622 580102
rect 589194 579922 589250 579978
rect 589318 579922 589374 579978
rect 589442 579922 589498 579978
rect 589566 579922 589622 579978
rect 27878 568294 27934 568350
rect 28002 568294 28058 568350
rect 27878 568170 27934 568226
rect 28002 568170 28058 568226
rect 27878 568046 27934 568102
rect 28002 568046 28058 568102
rect 27878 567922 27934 567978
rect 28002 567922 28058 567978
rect 58598 568294 58654 568350
rect 58722 568294 58778 568350
rect 58598 568170 58654 568226
rect 58722 568170 58778 568226
rect 58598 568046 58654 568102
rect 58722 568046 58778 568102
rect 58598 567922 58654 567978
rect 58722 567922 58778 567978
rect 89318 568294 89374 568350
rect 89442 568294 89498 568350
rect 89318 568170 89374 568226
rect 89442 568170 89498 568226
rect 89318 568046 89374 568102
rect 89442 568046 89498 568102
rect 89318 567922 89374 567978
rect 89442 567922 89498 567978
rect 120038 568294 120094 568350
rect 120162 568294 120218 568350
rect 120038 568170 120094 568226
rect 120162 568170 120218 568226
rect 120038 568046 120094 568102
rect 120162 568046 120218 568102
rect 120038 567922 120094 567978
rect 120162 567922 120218 567978
rect 150758 568294 150814 568350
rect 150882 568294 150938 568350
rect 150758 568170 150814 568226
rect 150882 568170 150938 568226
rect 150758 568046 150814 568102
rect 150882 568046 150938 568102
rect 150758 567922 150814 567978
rect 150882 567922 150938 567978
rect 181478 568294 181534 568350
rect 181602 568294 181658 568350
rect 181478 568170 181534 568226
rect 181602 568170 181658 568226
rect 181478 568046 181534 568102
rect 181602 568046 181658 568102
rect 181478 567922 181534 567978
rect 181602 567922 181658 567978
rect 212198 568294 212254 568350
rect 212322 568294 212378 568350
rect 212198 568170 212254 568226
rect 212322 568170 212378 568226
rect 212198 568046 212254 568102
rect 212322 568046 212378 568102
rect 212198 567922 212254 567978
rect 212322 567922 212378 567978
rect 242918 568294 242974 568350
rect 243042 568294 243098 568350
rect 242918 568170 242974 568226
rect 243042 568170 243098 568226
rect 242918 568046 242974 568102
rect 243042 568046 243098 568102
rect 242918 567922 242974 567978
rect 243042 567922 243098 567978
rect 273638 568294 273694 568350
rect 273762 568294 273818 568350
rect 273638 568170 273694 568226
rect 273762 568170 273818 568226
rect 273638 568046 273694 568102
rect 273762 568046 273818 568102
rect 273638 567922 273694 567978
rect 273762 567922 273818 567978
rect 304358 568294 304414 568350
rect 304482 568294 304538 568350
rect 304358 568170 304414 568226
rect 304482 568170 304538 568226
rect 304358 568046 304414 568102
rect 304482 568046 304538 568102
rect 304358 567922 304414 567978
rect 304482 567922 304538 567978
rect 335078 568294 335134 568350
rect 335202 568294 335258 568350
rect 335078 568170 335134 568226
rect 335202 568170 335258 568226
rect 335078 568046 335134 568102
rect 335202 568046 335258 568102
rect 335078 567922 335134 567978
rect 335202 567922 335258 567978
rect 365798 568294 365854 568350
rect 365922 568294 365978 568350
rect 365798 568170 365854 568226
rect 365922 568170 365978 568226
rect 365798 568046 365854 568102
rect 365922 568046 365978 568102
rect 365798 567922 365854 567978
rect 365922 567922 365978 567978
rect 396518 568294 396574 568350
rect 396642 568294 396698 568350
rect 396518 568170 396574 568226
rect 396642 568170 396698 568226
rect 396518 568046 396574 568102
rect 396642 568046 396698 568102
rect 396518 567922 396574 567978
rect 396642 567922 396698 567978
rect 427238 568294 427294 568350
rect 427362 568294 427418 568350
rect 427238 568170 427294 568226
rect 427362 568170 427418 568226
rect 427238 568046 427294 568102
rect 427362 568046 427418 568102
rect 427238 567922 427294 567978
rect 427362 567922 427418 567978
rect 457958 568294 458014 568350
rect 458082 568294 458138 568350
rect 457958 568170 458014 568226
rect 458082 568170 458138 568226
rect 457958 568046 458014 568102
rect 458082 568046 458138 568102
rect 457958 567922 458014 567978
rect 458082 567922 458138 567978
rect 488678 568294 488734 568350
rect 488802 568294 488858 568350
rect 488678 568170 488734 568226
rect 488802 568170 488858 568226
rect 488678 568046 488734 568102
rect 488802 568046 488858 568102
rect 488678 567922 488734 567978
rect 488802 567922 488858 567978
rect 519398 568294 519454 568350
rect 519522 568294 519578 568350
rect 519398 568170 519454 568226
rect 519522 568170 519578 568226
rect 519398 568046 519454 568102
rect 519522 568046 519578 568102
rect 519398 567922 519454 567978
rect 519522 567922 519578 567978
rect 550118 568294 550174 568350
rect 550242 568294 550298 568350
rect 550118 568170 550174 568226
rect 550242 568170 550298 568226
rect 550118 568046 550174 568102
rect 550242 568046 550298 568102
rect 550118 567922 550174 567978
rect 550242 567922 550298 567978
rect 5514 562294 5570 562350
rect 5638 562294 5694 562350
rect 5762 562294 5818 562350
rect 5886 562294 5942 562350
rect 5514 562170 5570 562226
rect 5638 562170 5694 562226
rect 5762 562170 5818 562226
rect 5886 562170 5942 562226
rect 5514 562046 5570 562102
rect 5638 562046 5694 562102
rect 5762 562046 5818 562102
rect 5886 562046 5942 562102
rect 5514 561922 5570 561978
rect 5638 561922 5694 561978
rect 5762 561922 5818 561978
rect 5886 561922 5942 561978
rect -860 544294 -804 544350
rect -736 544294 -680 544350
rect -612 544294 -556 544350
rect -488 544294 -432 544350
rect -860 544170 -804 544226
rect -736 544170 -680 544226
rect -612 544170 -556 544226
rect -488 544170 -432 544226
rect -860 544046 -804 544102
rect -736 544046 -680 544102
rect -612 544046 -556 544102
rect -488 544046 -432 544102
rect -860 543922 -804 543978
rect -736 543922 -680 543978
rect -612 543922 -556 543978
rect -488 543922 -432 543978
rect -860 526294 -804 526350
rect -736 526294 -680 526350
rect -612 526294 -556 526350
rect -488 526294 -432 526350
rect -860 526170 -804 526226
rect -736 526170 -680 526226
rect -612 526170 -556 526226
rect -488 526170 -432 526226
rect -860 526046 -804 526102
rect -736 526046 -680 526102
rect -612 526046 -556 526102
rect -488 526046 -432 526102
rect -860 525922 -804 525978
rect -736 525922 -680 525978
rect -612 525922 -556 525978
rect -488 525922 -432 525978
rect 12518 562294 12574 562350
rect 12642 562294 12698 562350
rect 12518 562170 12574 562226
rect 12642 562170 12698 562226
rect 12518 562046 12574 562102
rect 12642 562046 12698 562102
rect 12518 561922 12574 561978
rect 12642 561922 12698 561978
rect 43238 562294 43294 562350
rect 43362 562294 43418 562350
rect 43238 562170 43294 562226
rect 43362 562170 43418 562226
rect 43238 562046 43294 562102
rect 43362 562046 43418 562102
rect 43238 561922 43294 561978
rect 43362 561922 43418 561978
rect 73958 562294 74014 562350
rect 74082 562294 74138 562350
rect 73958 562170 74014 562226
rect 74082 562170 74138 562226
rect 73958 562046 74014 562102
rect 74082 562046 74138 562102
rect 73958 561922 74014 561978
rect 74082 561922 74138 561978
rect 104678 562294 104734 562350
rect 104802 562294 104858 562350
rect 104678 562170 104734 562226
rect 104802 562170 104858 562226
rect 104678 562046 104734 562102
rect 104802 562046 104858 562102
rect 104678 561922 104734 561978
rect 104802 561922 104858 561978
rect 135398 562294 135454 562350
rect 135522 562294 135578 562350
rect 135398 562170 135454 562226
rect 135522 562170 135578 562226
rect 135398 562046 135454 562102
rect 135522 562046 135578 562102
rect 135398 561922 135454 561978
rect 135522 561922 135578 561978
rect 166118 562294 166174 562350
rect 166242 562294 166298 562350
rect 166118 562170 166174 562226
rect 166242 562170 166298 562226
rect 166118 562046 166174 562102
rect 166242 562046 166298 562102
rect 166118 561922 166174 561978
rect 166242 561922 166298 561978
rect 196838 562294 196894 562350
rect 196962 562294 197018 562350
rect 196838 562170 196894 562226
rect 196962 562170 197018 562226
rect 196838 562046 196894 562102
rect 196962 562046 197018 562102
rect 196838 561922 196894 561978
rect 196962 561922 197018 561978
rect 227558 562294 227614 562350
rect 227682 562294 227738 562350
rect 227558 562170 227614 562226
rect 227682 562170 227738 562226
rect 227558 562046 227614 562102
rect 227682 562046 227738 562102
rect 227558 561922 227614 561978
rect 227682 561922 227738 561978
rect 258278 562294 258334 562350
rect 258402 562294 258458 562350
rect 258278 562170 258334 562226
rect 258402 562170 258458 562226
rect 258278 562046 258334 562102
rect 258402 562046 258458 562102
rect 258278 561922 258334 561978
rect 258402 561922 258458 561978
rect 288998 562294 289054 562350
rect 289122 562294 289178 562350
rect 288998 562170 289054 562226
rect 289122 562170 289178 562226
rect 288998 562046 289054 562102
rect 289122 562046 289178 562102
rect 288998 561922 289054 561978
rect 289122 561922 289178 561978
rect 319718 562294 319774 562350
rect 319842 562294 319898 562350
rect 319718 562170 319774 562226
rect 319842 562170 319898 562226
rect 319718 562046 319774 562102
rect 319842 562046 319898 562102
rect 319718 561922 319774 561978
rect 319842 561922 319898 561978
rect 350438 562294 350494 562350
rect 350562 562294 350618 562350
rect 350438 562170 350494 562226
rect 350562 562170 350618 562226
rect 350438 562046 350494 562102
rect 350562 562046 350618 562102
rect 350438 561922 350494 561978
rect 350562 561922 350618 561978
rect 381158 562294 381214 562350
rect 381282 562294 381338 562350
rect 381158 562170 381214 562226
rect 381282 562170 381338 562226
rect 381158 562046 381214 562102
rect 381282 562046 381338 562102
rect 381158 561922 381214 561978
rect 381282 561922 381338 561978
rect 411878 562294 411934 562350
rect 412002 562294 412058 562350
rect 411878 562170 411934 562226
rect 412002 562170 412058 562226
rect 411878 562046 411934 562102
rect 412002 562046 412058 562102
rect 411878 561922 411934 561978
rect 412002 561922 412058 561978
rect 442598 562294 442654 562350
rect 442722 562294 442778 562350
rect 442598 562170 442654 562226
rect 442722 562170 442778 562226
rect 442598 562046 442654 562102
rect 442722 562046 442778 562102
rect 442598 561922 442654 561978
rect 442722 561922 442778 561978
rect 473318 562294 473374 562350
rect 473442 562294 473498 562350
rect 473318 562170 473374 562226
rect 473442 562170 473498 562226
rect 473318 562046 473374 562102
rect 473442 562046 473498 562102
rect 473318 561922 473374 561978
rect 473442 561922 473498 561978
rect 504038 562294 504094 562350
rect 504162 562294 504218 562350
rect 504038 562170 504094 562226
rect 504162 562170 504218 562226
rect 504038 562046 504094 562102
rect 504162 562046 504218 562102
rect 504038 561922 504094 561978
rect 504162 561922 504218 561978
rect 534758 562294 534814 562350
rect 534882 562294 534938 562350
rect 534758 562170 534814 562226
rect 534882 562170 534938 562226
rect 534758 562046 534814 562102
rect 534882 562046 534938 562102
rect 534758 561922 534814 561978
rect 534882 561922 534938 561978
rect 565478 562294 565534 562350
rect 565602 562294 565658 562350
rect 565478 562170 565534 562226
rect 565602 562170 565658 562226
rect 597456 598116 597512 598172
rect 597580 598116 597636 598172
rect 597704 598116 597760 598172
rect 597828 598116 597884 598172
rect 597456 597992 597512 598048
rect 597580 597992 597636 598048
rect 597704 597992 597760 598048
rect 597828 597992 597884 598048
rect 597456 597868 597512 597924
rect 597580 597868 597636 597924
rect 597704 597868 597760 597924
rect 597828 597868 597884 597924
rect 597456 597744 597512 597800
rect 597580 597744 597636 597800
rect 597704 597744 597760 597800
rect 597828 597744 597884 597800
rect 592914 586294 592970 586350
rect 593038 586294 593094 586350
rect 593162 586294 593218 586350
rect 593286 586294 593342 586350
rect 592914 586170 592970 586226
rect 593038 586170 593094 586226
rect 593162 586170 593218 586226
rect 593286 586170 593342 586226
rect 592914 586046 592970 586102
rect 593038 586046 593094 586102
rect 593162 586046 593218 586102
rect 593286 586046 593342 586102
rect 592914 585922 592970 585978
rect 593038 585922 593094 585978
rect 593162 585922 593218 585978
rect 593286 585922 593342 585978
rect 592914 568294 592970 568350
rect 593038 568294 593094 568350
rect 593162 568294 593218 568350
rect 593286 568294 593342 568350
rect 592914 568170 592970 568226
rect 593038 568170 593094 568226
rect 593162 568170 593218 568226
rect 593286 568170 593342 568226
rect 592914 568046 592970 568102
rect 593038 568046 593094 568102
rect 593162 568046 593218 568102
rect 593286 568046 593342 568102
rect 592914 567922 592970 567978
rect 593038 567922 593094 567978
rect 593162 567922 593218 567978
rect 593286 567922 593342 567978
rect 589194 562294 589250 562350
rect 589318 562294 589374 562350
rect 589442 562294 589498 562350
rect 589566 562294 589622 562350
rect 565478 562046 565534 562102
rect 565602 562046 565658 562102
rect 565478 561922 565534 561978
rect 565602 561922 565658 561978
rect 5514 544294 5570 544350
rect 5638 544294 5694 544350
rect 5762 544294 5818 544350
rect 5886 544294 5942 544350
rect 5514 544170 5570 544226
rect 5638 544170 5694 544226
rect 5762 544170 5818 544226
rect 5886 544170 5942 544226
rect 5514 544046 5570 544102
rect 5638 544046 5694 544102
rect 5762 544046 5818 544102
rect 5886 544046 5942 544102
rect 589194 562170 589250 562226
rect 589318 562170 589374 562226
rect 589442 562170 589498 562226
rect 589566 562170 589622 562226
rect 589194 562046 589250 562102
rect 589318 562046 589374 562102
rect 589442 562046 589498 562102
rect 589566 562046 589622 562102
rect 589194 561922 589250 561978
rect 589318 561922 589374 561978
rect 589442 561922 589498 561978
rect 589566 561922 589622 561978
rect 27878 550294 27934 550350
rect 28002 550294 28058 550350
rect 27878 550170 27934 550226
rect 28002 550170 28058 550226
rect 27878 550046 27934 550102
rect 28002 550046 28058 550102
rect 27878 549922 27934 549978
rect 28002 549922 28058 549978
rect 58598 550294 58654 550350
rect 58722 550294 58778 550350
rect 58598 550170 58654 550226
rect 58722 550170 58778 550226
rect 58598 550046 58654 550102
rect 58722 550046 58778 550102
rect 58598 549922 58654 549978
rect 58722 549922 58778 549978
rect 89318 550294 89374 550350
rect 89442 550294 89498 550350
rect 89318 550170 89374 550226
rect 89442 550170 89498 550226
rect 89318 550046 89374 550102
rect 89442 550046 89498 550102
rect 89318 549922 89374 549978
rect 89442 549922 89498 549978
rect 120038 550294 120094 550350
rect 120162 550294 120218 550350
rect 120038 550170 120094 550226
rect 120162 550170 120218 550226
rect 120038 550046 120094 550102
rect 120162 550046 120218 550102
rect 120038 549922 120094 549978
rect 120162 549922 120218 549978
rect 150758 550294 150814 550350
rect 150882 550294 150938 550350
rect 150758 550170 150814 550226
rect 150882 550170 150938 550226
rect 150758 550046 150814 550102
rect 150882 550046 150938 550102
rect 150758 549922 150814 549978
rect 150882 549922 150938 549978
rect 181478 550294 181534 550350
rect 181602 550294 181658 550350
rect 181478 550170 181534 550226
rect 181602 550170 181658 550226
rect 181478 550046 181534 550102
rect 181602 550046 181658 550102
rect 181478 549922 181534 549978
rect 181602 549922 181658 549978
rect 212198 550294 212254 550350
rect 212322 550294 212378 550350
rect 212198 550170 212254 550226
rect 212322 550170 212378 550226
rect 212198 550046 212254 550102
rect 212322 550046 212378 550102
rect 212198 549922 212254 549978
rect 212322 549922 212378 549978
rect 242918 550294 242974 550350
rect 243042 550294 243098 550350
rect 242918 550170 242974 550226
rect 243042 550170 243098 550226
rect 242918 550046 242974 550102
rect 243042 550046 243098 550102
rect 242918 549922 242974 549978
rect 243042 549922 243098 549978
rect 273638 550294 273694 550350
rect 273762 550294 273818 550350
rect 273638 550170 273694 550226
rect 273762 550170 273818 550226
rect 273638 550046 273694 550102
rect 273762 550046 273818 550102
rect 273638 549922 273694 549978
rect 273762 549922 273818 549978
rect 304358 550294 304414 550350
rect 304482 550294 304538 550350
rect 304358 550170 304414 550226
rect 304482 550170 304538 550226
rect 304358 550046 304414 550102
rect 304482 550046 304538 550102
rect 304358 549922 304414 549978
rect 304482 549922 304538 549978
rect 335078 550294 335134 550350
rect 335202 550294 335258 550350
rect 335078 550170 335134 550226
rect 335202 550170 335258 550226
rect 335078 550046 335134 550102
rect 335202 550046 335258 550102
rect 335078 549922 335134 549978
rect 335202 549922 335258 549978
rect 365798 550294 365854 550350
rect 365922 550294 365978 550350
rect 365798 550170 365854 550226
rect 365922 550170 365978 550226
rect 365798 550046 365854 550102
rect 365922 550046 365978 550102
rect 365798 549922 365854 549978
rect 365922 549922 365978 549978
rect 396518 550294 396574 550350
rect 396642 550294 396698 550350
rect 396518 550170 396574 550226
rect 396642 550170 396698 550226
rect 396518 550046 396574 550102
rect 396642 550046 396698 550102
rect 396518 549922 396574 549978
rect 396642 549922 396698 549978
rect 427238 550294 427294 550350
rect 427362 550294 427418 550350
rect 427238 550170 427294 550226
rect 427362 550170 427418 550226
rect 427238 550046 427294 550102
rect 427362 550046 427418 550102
rect 427238 549922 427294 549978
rect 427362 549922 427418 549978
rect 457958 550294 458014 550350
rect 458082 550294 458138 550350
rect 457958 550170 458014 550226
rect 458082 550170 458138 550226
rect 457958 550046 458014 550102
rect 458082 550046 458138 550102
rect 457958 549922 458014 549978
rect 458082 549922 458138 549978
rect 488678 550294 488734 550350
rect 488802 550294 488858 550350
rect 488678 550170 488734 550226
rect 488802 550170 488858 550226
rect 488678 550046 488734 550102
rect 488802 550046 488858 550102
rect 488678 549922 488734 549978
rect 488802 549922 488858 549978
rect 519398 550294 519454 550350
rect 519522 550294 519578 550350
rect 519398 550170 519454 550226
rect 519522 550170 519578 550226
rect 519398 550046 519454 550102
rect 519522 550046 519578 550102
rect 519398 549922 519454 549978
rect 519522 549922 519578 549978
rect 550118 550294 550174 550350
rect 550242 550294 550298 550350
rect 550118 550170 550174 550226
rect 550242 550170 550298 550226
rect 550118 550046 550174 550102
rect 550242 550046 550298 550102
rect 550118 549922 550174 549978
rect 550242 549922 550298 549978
rect 12518 544294 12574 544350
rect 12642 544294 12698 544350
rect 12518 544170 12574 544226
rect 12642 544170 12698 544226
rect 12518 544046 12574 544102
rect 12642 544046 12698 544102
rect 5514 543922 5570 543978
rect 5638 543922 5694 543978
rect 5762 543922 5818 543978
rect 5886 543922 5942 543978
rect 12518 543922 12574 543978
rect 12642 543922 12698 543978
rect 43238 544294 43294 544350
rect 43362 544294 43418 544350
rect 43238 544170 43294 544226
rect 43362 544170 43418 544226
rect 43238 544046 43294 544102
rect 43362 544046 43418 544102
rect 43238 543922 43294 543978
rect 43362 543922 43418 543978
rect 73958 544294 74014 544350
rect 74082 544294 74138 544350
rect 73958 544170 74014 544226
rect 74082 544170 74138 544226
rect 73958 544046 74014 544102
rect 74082 544046 74138 544102
rect 73958 543922 74014 543978
rect 74082 543922 74138 543978
rect 104678 544294 104734 544350
rect 104802 544294 104858 544350
rect 104678 544170 104734 544226
rect 104802 544170 104858 544226
rect 104678 544046 104734 544102
rect 104802 544046 104858 544102
rect 104678 543922 104734 543978
rect 104802 543922 104858 543978
rect 135398 544294 135454 544350
rect 135522 544294 135578 544350
rect 135398 544170 135454 544226
rect 135522 544170 135578 544226
rect 135398 544046 135454 544102
rect 135522 544046 135578 544102
rect 135398 543922 135454 543978
rect 135522 543922 135578 543978
rect 166118 544294 166174 544350
rect 166242 544294 166298 544350
rect 166118 544170 166174 544226
rect 166242 544170 166298 544226
rect 166118 544046 166174 544102
rect 166242 544046 166298 544102
rect 166118 543922 166174 543978
rect 166242 543922 166298 543978
rect 196838 544294 196894 544350
rect 196962 544294 197018 544350
rect 196838 544170 196894 544226
rect 196962 544170 197018 544226
rect 196838 544046 196894 544102
rect 196962 544046 197018 544102
rect 196838 543922 196894 543978
rect 196962 543922 197018 543978
rect 227558 544294 227614 544350
rect 227682 544294 227738 544350
rect 227558 544170 227614 544226
rect 227682 544170 227738 544226
rect 227558 544046 227614 544102
rect 227682 544046 227738 544102
rect 227558 543922 227614 543978
rect 227682 543922 227738 543978
rect 258278 544294 258334 544350
rect 258402 544294 258458 544350
rect 258278 544170 258334 544226
rect 258402 544170 258458 544226
rect 258278 544046 258334 544102
rect 258402 544046 258458 544102
rect 258278 543922 258334 543978
rect 258402 543922 258458 543978
rect 288998 544294 289054 544350
rect 289122 544294 289178 544350
rect 288998 544170 289054 544226
rect 289122 544170 289178 544226
rect 288998 544046 289054 544102
rect 289122 544046 289178 544102
rect 288998 543922 289054 543978
rect 289122 543922 289178 543978
rect 319718 544294 319774 544350
rect 319842 544294 319898 544350
rect 319718 544170 319774 544226
rect 319842 544170 319898 544226
rect 319718 544046 319774 544102
rect 319842 544046 319898 544102
rect 319718 543922 319774 543978
rect 319842 543922 319898 543978
rect 350438 544294 350494 544350
rect 350562 544294 350618 544350
rect 350438 544170 350494 544226
rect 350562 544170 350618 544226
rect 350438 544046 350494 544102
rect 350562 544046 350618 544102
rect 350438 543922 350494 543978
rect 350562 543922 350618 543978
rect 381158 544294 381214 544350
rect 381282 544294 381338 544350
rect 381158 544170 381214 544226
rect 381282 544170 381338 544226
rect 381158 544046 381214 544102
rect 381282 544046 381338 544102
rect 381158 543922 381214 543978
rect 381282 543922 381338 543978
rect 411878 544294 411934 544350
rect 412002 544294 412058 544350
rect 411878 544170 411934 544226
rect 412002 544170 412058 544226
rect 411878 544046 411934 544102
rect 412002 544046 412058 544102
rect 411878 543922 411934 543978
rect 412002 543922 412058 543978
rect 442598 544294 442654 544350
rect 442722 544294 442778 544350
rect 442598 544170 442654 544226
rect 442722 544170 442778 544226
rect 442598 544046 442654 544102
rect 442722 544046 442778 544102
rect 442598 543922 442654 543978
rect 442722 543922 442778 543978
rect 473318 544294 473374 544350
rect 473442 544294 473498 544350
rect 473318 544170 473374 544226
rect 473442 544170 473498 544226
rect 473318 544046 473374 544102
rect 473442 544046 473498 544102
rect 473318 543922 473374 543978
rect 473442 543922 473498 543978
rect 504038 544294 504094 544350
rect 504162 544294 504218 544350
rect 504038 544170 504094 544226
rect 504162 544170 504218 544226
rect 504038 544046 504094 544102
rect 504162 544046 504218 544102
rect 504038 543922 504094 543978
rect 504162 543922 504218 543978
rect 534758 544294 534814 544350
rect 534882 544294 534938 544350
rect 534758 544170 534814 544226
rect 534882 544170 534938 544226
rect 534758 544046 534814 544102
rect 534882 544046 534938 544102
rect 534758 543922 534814 543978
rect 534882 543922 534938 543978
rect 565478 544294 565534 544350
rect 565602 544294 565658 544350
rect 565478 544170 565534 544226
rect 565602 544170 565658 544226
rect 565478 544046 565534 544102
rect 565602 544046 565658 544102
rect 565478 543922 565534 543978
rect 565602 543922 565658 543978
rect 592914 550294 592970 550350
rect 593038 550294 593094 550350
rect 593162 550294 593218 550350
rect 593286 550294 593342 550350
rect 592914 550170 592970 550226
rect 593038 550170 593094 550226
rect 593162 550170 593218 550226
rect 593286 550170 593342 550226
rect 592914 550046 592970 550102
rect 593038 550046 593094 550102
rect 593162 550046 593218 550102
rect 593286 550046 593342 550102
rect 592914 549922 592970 549978
rect 593038 549922 593094 549978
rect 593162 549922 593218 549978
rect 593286 549922 593342 549978
rect 589194 544294 589250 544350
rect 589318 544294 589374 544350
rect 589442 544294 589498 544350
rect 589566 544294 589622 544350
rect 589194 544170 589250 544226
rect 589318 544170 589374 544226
rect 589442 544170 589498 544226
rect 589566 544170 589622 544226
rect 589194 544046 589250 544102
rect 589318 544046 589374 544102
rect 589442 544046 589498 544102
rect 589566 544046 589622 544102
rect 589194 543922 589250 543978
rect 589318 543922 589374 543978
rect 589442 543922 589498 543978
rect 589566 543922 589622 543978
rect 27878 532294 27934 532350
rect 28002 532294 28058 532350
rect 27878 532170 27934 532226
rect 28002 532170 28058 532226
rect 27878 532046 27934 532102
rect 28002 532046 28058 532102
rect 27878 531922 27934 531978
rect 28002 531922 28058 531978
rect 58598 532294 58654 532350
rect 58722 532294 58778 532350
rect 58598 532170 58654 532226
rect 58722 532170 58778 532226
rect 58598 532046 58654 532102
rect 58722 532046 58778 532102
rect 58598 531922 58654 531978
rect 58722 531922 58778 531978
rect 89318 532294 89374 532350
rect 89442 532294 89498 532350
rect 89318 532170 89374 532226
rect 89442 532170 89498 532226
rect 89318 532046 89374 532102
rect 89442 532046 89498 532102
rect 89318 531922 89374 531978
rect 89442 531922 89498 531978
rect 120038 532294 120094 532350
rect 120162 532294 120218 532350
rect 120038 532170 120094 532226
rect 120162 532170 120218 532226
rect 120038 532046 120094 532102
rect 120162 532046 120218 532102
rect 120038 531922 120094 531978
rect 120162 531922 120218 531978
rect 150758 532294 150814 532350
rect 150882 532294 150938 532350
rect 150758 532170 150814 532226
rect 150882 532170 150938 532226
rect 150758 532046 150814 532102
rect 150882 532046 150938 532102
rect 150758 531922 150814 531978
rect 150882 531922 150938 531978
rect 181478 532294 181534 532350
rect 181602 532294 181658 532350
rect 181478 532170 181534 532226
rect 181602 532170 181658 532226
rect 181478 532046 181534 532102
rect 181602 532046 181658 532102
rect 181478 531922 181534 531978
rect 181602 531922 181658 531978
rect 212198 532294 212254 532350
rect 212322 532294 212378 532350
rect 212198 532170 212254 532226
rect 212322 532170 212378 532226
rect 212198 532046 212254 532102
rect 212322 532046 212378 532102
rect 212198 531922 212254 531978
rect 212322 531922 212378 531978
rect 242918 532294 242974 532350
rect 243042 532294 243098 532350
rect 242918 532170 242974 532226
rect 243042 532170 243098 532226
rect 242918 532046 242974 532102
rect 243042 532046 243098 532102
rect 242918 531922 242974 531978
rect 243042 531922 243098 531978
rect 273638 532294 273694 532350
rect 273762 532294 273818 532350
rect 273638 532170 273694 532226
rect 273762 532170 273818 532226
rect 273638 532046 273694 532102
rect 273762 532046 273818 532102
rect 273638 531922 273694 531978
rect 273762 531922 273818 531978
rect 304358 532294 304414 532350
rect 304482 532294 304538 532350
rect 304358 532170 304414 532226
rect 304482 532170 304538 532226
rect 304358 532046 304414 532102
rect 304482 532046 304538 532102
rect 304358 531922 304414 531978
rect 304482 531922 304538 531978
rect 335078 532294 335134 532350
rect 335202 532294 335258 532350
rect 335078 532170 335134 532226
rect 335202 532170 335258 532226
rect 335078 532046 335134 532102
rect 335202 532046 335258 532102
rect 335078 531922 335134 531978
rect 335202 531922 335258 531978
rect 365798 532294 365854 532350
rect 365922 532294 365978 532350
rect 365798 532170 365854 532226
rect 365922 532170 365978 532226
rect 365798 532046 365854 532102
rect 365922 532046 365978 532102
rect 365798 531922 365854 531978
rect 365922 531922 365978 531978
rect 396518 532294 396574 532350
rect 396642 532294 396698 532350
rect 396518 532170 396574 532226
rect 396642 532170 396698 532226
rect 396518 532046 396574 532102
rect 396642 532046 396698 532102
rect 396518 531922 396574 531978
rect 396642 531922 396698 531978
rect 427238 532294 427294 532350
rect 427362 532294 427418 532350
rect 427238 532170 427294 532226
rect 427362 532170 427418 532226
rect 427238 532046 427294 532102
rect 427362 532046 427418 532102
rect 427238 531922 427294 531978
rect 427362 531922 427418 531978
rect 457958 532294 458014 532350
rect 458082 532294 458138 532350
rect 457958 532170 458014 532226
rect 458082 532170 458138 532226
rect 457958 532046 458014 532102
rect 458082 532046 458138 532102
rect 457958 531922 458014 531978
rect 458082 531922 458138 531978
rect 488678 532294 488734 532350
rect 488802 532294 488858 532350
rect 488678 532170 488734 532226
rect 488802 532170 488858 532226
rect 488678 532046 488734 532102
rect 488802 532046 488858 532102
rect 488678 531922 488734 531978
rect 488802 531922 488858 531978
rect 519398 532294 519454 532350
rect 519522 532294 519578 532350
rect 519398 532170 519454 532226
rect 519522 532170 519578 532226
rect 519398 532046 519454 532102
rect 519522 532046 519578 532102
rect 519398 531922 519454 531978
rect 519522 531922 519578 531978
rect 550118 532294 550174 532350
rect 550242 532294 550298 532350
rect 550118 532170 550174 532226
rect 550242 532170 550298 532226
rect 550118 532046 550174 532102
rect 550242 532046 550298 532102
rect 550118 531922 550174 531978
rect 550242 531922 550298 531978
rect 5514 526294 5570 526350
rect 5638 526294 5694 526350
rect 5762 526294 5818 526350
rect 5886 526294 5942 526350
rect 5514 526170 5570 526226
rect 5638 526170 5694 526226
rect 5762 526170 5818 526226
rect 5886 526170 5942 526226
rect 5514 526046 5570 526102
rect 5638 526046 5694 526102
rect 5762 526046 5818 526102
rect 5886 526046 5942 526102
rect 5514 525922 5570 525978
rect 5638 525922 5694 525978
rect 5762 525922 5818 525978
rect 5886 525922 5942 525978
rect -860 508294 -804 508350
rect -736 508294 -680 508350
rect -612 508294 -556 508350
rect -488 508294 -432 508350
rect -860 508170 -804 508226
rect -736 508170 -680 508226
rect -612 508170 -556 508226
rect -488 508170 -432 508226
rect -860 508046 -804 508102
rect -736 508046 -680 508102
rect -612 508046 -556 508102
rect -488 508046 -432 508102
rect -860 507922 -804 507978
rect -736 507922 -680 507978
rect -612 507922 -556 507978
rect -488 507922 -432 507978
rect 12518 526294 12574 526350
rect 12642 526294 12698 526350
rect 12518 526170 12574 526226
rect 12642 526170 12698 526226
rect 12518 526046 12574 526102
rect 12642 526046 12698 526102
rect 12518 525922 12574 525978
rect 12642 525922 12698 525978
rect 43238 526294 43294 526350
rect 43362 526294 43418 526350
rect 43238 526170 43294 526226
rect 43362 526170 43418 526226
rect 43238 526046 43294 526102
rect 43362 526046 43418 526102
rect 43238 525922 43294 525978
rect 43362 525922 43418 525978
rect 73958 526294 74014 526350
rect 74082 526294 74138 526350
rect 73958 526170 74014 526226
rect 74082 526170 74138 526226
rect 73958 526046 74014 526102
rect 74082 526046 74138 526102
rect 73958 525922 74014 525978
rect 74082 525922 74138 525978
rect 104678 526294 104734 526350
rect 104802 526294 104858 526350
rect 104678 526170 104734 526226
rect 104802 526170 104858 526226
rect 104678 526046 104734 526102
rect 104802 526046 104858 526102
rect 104678 525922 104734 525978
rect 104802 525922 104858 525978
rect 135398 526294 135454 526350
rect 135522 526294 135578 526350
rect 135398 526170 135454 526226
rect 135522 526170 135578 526226
rect 135398 526046 135454 526102
rect 135522 526046 135578 526102
rect 135398 525922 135454 525978
rect 135522 525922 135578 525978
rect 166118 526294 166174 526350
rect 166242 526294 166298 526350
rect 166118 526170 166174 526226
rect 166242 526170 166298 526226
rect 166118 526046 166174 526102
rect 166242 526046 166298 526102
rect 166118 525922 166174 525978
rect 166242 525922 166298 525978
rect 196838 526294 196894 526350
rect 196962 526294 197018 526350
rect 196838 526170 196894 526226
rect 196962 526170 197018 526226
rect 196838 526046 196894 526102
rect 196962 526046 197018 526102
rect 196838 525922 196894 525978
rect 196962 525922 197018 525978
rect 227558 526294 227614 526350
rect 227682 526294 227738 526350
rect 227558 526170 227614 526226
rect 227682 526170 227738 526226
rect 227558 526046 227614 526102
rect 227682 526046 227738 526102
rect 227558 525922 227614 525978
rect 227682 525922 227738 525978
rect 258278 526294 258334 526350
rect 258402 526294 258458 526350
rect 258278 526170 258334 526226
rect 258402 526170 258458 526226
rect 258278 526046 258334 526102
rect 258402 526046 258458 526102
rect 258278 525922 258334 525978
rect 258402 525922 258458 525978
rect 288998 526294 289054 526350
rect 289122 526294 289178 526350
rect 288998 526170 289054 526226
rect 289122 526170 289178 526226
rect 288998 526046 289054 526102
rect 289122 526046 289178 526102
rect 288998 525922 289054 525978
rect 289122 525922 289178 525978
rect 319718 526294 319774 526350
rect 319842 526294 319898 526350
rect 319718 526170 319774 526226
rect 319842 526170 319898 526226
rect 319718 526046 319774 526102
rect 319842 526046 319898 526102
rect 319718 525922 319774 525978
rect 319842 525922 319898 525978
rect 350438 526294 350494 526350
rect 350562 526294 350618 526350
rect 350438 526170 350494 526226
rect 350562 526170 350618 526226
rect 350438 526046 350494 526102
rect 350562 526046 350618 526102
rect 350438 525922 350494 525978
rect 350562 525922 350618 525978
rect 381158 526294 381214 526350
rect 381282 526294 381338 526350
rect 381158 526170 381214 526226
rect 381282 526170 381338 526226
rect 381158 526046 381214 526102
rect 381282 526046 381338 526102
rect 381158 525922 381214 525978
rect 381282 525922 381338 525978
rect 411878 526294 411934 526350
rect 412002 526294 412058 526350
rect 411878 526170 411934 526226
rect 412002 526170 412058 526226
rect 411878 526046 411934 526102
rect 412002 526046 412058 526102
rect 411878 525922 411934 525978
rect 412002 525922 412058 525978
rect 442598 526294 442654 526350
rect 442722 526294 442778 526350
rect 442598 526170 442654 526226
rect 442722 526170 442778 526226
rect 442598 526046 442654 526102
rect 442722 526046 442778 526102
rect 442598 525922 442654 525978
rect 442722 525922 442778 525978
rect 473318 526294 473374 526350
rect 473442 526294 473498 526350
rect 473318 526170 473374 526226
rect 473442 526170 473498 526226
rect 473318 526046 473374 526102
rect 473442 526046 473498 526102
rect 473318 525922 473374 525978
rect 473442 525922 473498 525978
rect 504038 526294 504094 526350
rect 504162 526294 504218 526350
rect 504038 526170 504094 526226
rect 504162 526170 504218 526226
rect 504038 526046 504094 526102
rect 504162 526046 504218 526102
rect 504038 525922 504094 525978
rect 504162 525922 504218 525978
rect 534758 526294 534814 526350
rect 534882 526294 534938 526350
rect 534758 526170 534814 526226
rect 534882 526170 534938 526226
rect 534758 526046 534814 526102
rect 534882 526046 534938 526102
rect 534758 525922 534814 525978
rect 534882 525922 534938 525978
rect 565478 526294 565534 526350
rect 565602 526294 565658 526350
rect 565478 526170 565534 526226
rect 565602 526170 565658 526226
rect 565478 526046 565534 526102
rect 565602 526046 565658 526102
rect 565478 525922 565534 525978
rect 565602 525922 565658 525978
rect 589194 526294 589250 526350
rect 589318 526294 589374 526350
rect 589442 526294 589498 526350
rect 589566 526294 589622 526350
rect 589194 526170 589250 526226
rect 589318 526170 589374 526226
rect 589442 526170 589498 526226
rect 589566 526170 589622 526226
rect 589194 526046 589250 526102
rect 589318 526046 589374 526102
rect 589442 526046 589498 526102
rect 589566 526046 589622 526102
rect 589194 525922 589250 525978
rect 589318 525922 589374 525978
rect 589442 525922 589498 525978
rect 589566 525922 589622 525978
rect 5514 508294 5570 508350
rect 5638 508294 5694 508350
rect 5762 508294 5818 508350
rect 5886 508294 5942 508350
rect 5514 508170 5570 508226
rect 5638 508170 5694 508226
rect 5762 508170 5818 508226
rect 5886 508170 5942 508226
rect 5514 508046 5570 508102
rect 5638 508046 5694 508102
rect 5762 508046 5818 508102
rect 5886 508046 5942 508102
rect 5514 507922 5570 507978
rect 5638 507922 5694 507978
rect 5762 507922 5818 507978
rect 5886 507922 5942 507978
rect -860 490294 -804 490350
rect -736 490294 -680 490350
rect -612 490294 -556 490350
rect -488 490294 -432 490350
rect -860 490170 -804 490226
rect -736 490170 -680 490226
rect -612 490170 -556 490226
rect -488 490170 -432 490226
rect -860 490046 -804 490102
rect -736 490046 -680 490102
rect -612 490046 -556 490102
rect -488 490046 -432 490102
rect -860 489922 -804 489978
rect -736 489922 -680 489978
rect -612 489922 -556 489978
rect -488 489922 -432 489978
rect 27878 514294 27934 514350
rect 28002 514294 28058 514350
rect 27878 514170 27934 514226
rect 28002 514170 28058 514226
rect 27878 514046 27934 514102
rect 28002 514046 28058 514102
rect 27878 513922 27934 513978
rect 28002 513922 28058 513978
rect 58598 514294 58654 514350
rect 58722 514294 58778 514350
rect 58598 514170 58654 514226
rect 58722 514170 58778 514226
rect 58598 514046 58654 514102
rect 58722 514046 58778 514102
rect 58598 513922 58654 513978
rect 58722 513922 58778 513978
rect 89318 514294 89374 514350
rect 89442 514294 89498 514350
rect 89318 514170 89374 514226
rect 89442 514170 89498 514226
rect 89318 514046 89374 514102
rect 89442 514046 89498 514102
rect 89318 513922 89374 513978
rect 89442 513922 89498 513978
rect 120038 514294 120094 514350
rect 120162 514294 120218 514350
rect 120038 514170 120094 514226
rect 120162 514170 120218 514226
rect 120038 514046 120094 514102
rect 120162 514046 120218 514102
rect 120038 513922 120094 513978
rect 120162 513922 120218 513978
rect 150758 514294 150814 514350
rect 150882 514294 150938 514350
rect 150758 514170 150814 514226
rect 150882 514170 150938 514226
rect 150758 514046 150814 514102
rect 150882 514046 150938 514102
rect 150758 513922 150814 513978
rect 150882 513922 150938 513978
rect 181478 514294 181534 514350
rect 181602 514294 181658 514350
rect 181478 514170 181534 514226
rect 181602 514170 181658 514226
rect 181478 514046 181534 514102
rect 181602 514046 181658 514102
rect 181478 513922 181534 513978
rect 181602 513922 181658 513978
rect 212198 514294 212254 514350
rect 212322 514294 212378 514350
rect 212198 514170 212254 514226
rect 212322 514170 212378 514226
rect 212198 514046 212254 514102
rect 212322 514046 212378 514102
rect 212198 513922 212254 513978
rect 212322 513922 212378 513978
rect 242918 514294 242974 514350
rect 243042 514294 243098 514350
rect 242918 514170 242974 514226
rect 243042 514170 243098 514226
rect 242918 514046 242974 514102
rect 243042 514046 243098 514102
rect 242918 513922 242974 513978
rect 243042 513922 243098 513978
rect 273638 514294 273694 514350
rect 273762 514294 273818 514350
rect 273638 514170 273694 514226
rect 273762 514170 273818 514226
rect 273638 514046 273694 514102
rect 273762 514046 273818 514102
rect 273638 513922 273694 513978
rect 273762 513922 273818 513978
rect 304358 514294 304414 514350
rect 304482 514294 304538 514350
rect 304358 514170 304414 514226
rect 304482 514170 304538 514226
rect 304358 514046 304414 514102
rect 304482 514046 304538 514102
rect 304358 513922 304414 513978
rect 304482 513922 304538 513978
rect 335078 514294 335134 514350
rect 335202 514294 335258 514350
rect 335078 514170 335134 514226
rect 335202 514170 335258 514226
rect 335078 514046 335134 514102
rect 335202 514046 335258 514102
rect 335078 513922 335134 513978
rect 335202 513922 335258 513978
rect 365798 514294 365854 514350
rect 365922 514294 365978 514350
rect 365798 514170 365854 514226
rect 365922 514170 365978 514226
rect 365798 514046 365854 514102
rect 365922 514046 365978 514102
rect 365798 513922 365854 513978
rect 365922 513922 365978 513978
rect 396518 514294 396574 514350
rect 396642 514294 396698 514350
rect 396518 514170 396574 514226
rect 396642 514170 396698 514226
rect 396518 514046 396574 514102
rect 396642 514046 396698 514102
rect 396518 513922 396574 513978
rect 396642 513922 396698 513978
rect 427238 514294 427294 514350
rect 427362 514294 427418 514350
rect 427238 514170 427294 514226
rect 427362 514170 427418 514226
rect 427238 514046 427294 514102
rect 427362 514046 427418 514102
rect 427238 513922 427294 513978
rect 427362 513922 427418 513978
rect 457958 514294 458014 514350
rect 458082 514294 458138 514350
rect 457958 514170 458014 514226
rect 458082 514170 458138 514226
rect 457958 514046 458014 514102
rect 458082 514046 458138 514102
rect 457958 513922 458014 513978
rect 458082 513922 458138 513978
rect 488678 514294 488734 514350
rect 488802 514294 488858 514350
rect 488678 514170 488734 514226
rect 488802 514170 488858 514226
rect 488678 514046 488734 514102
rect 488802 514046 488858 514102
rect 488678 513922 488734 513978
rect 488802 513922 488858 513978
rect 519398 514294 519454 514350
rect 519522 514294 519578 514350
rect 519398 514170 519454 514226
rect 519522 514170 519578 514226
rect 519398 514046 519454 514102
rect 519522 514046 519578 514102
rect 519398 513922 519454 513978
rect 519522 513922 519578 513978
rect 550118 514294 550174 514350
rect 550242 514294 550298 514350
rect 550118 514170 550174 514226
rect 550242 514170 550298 514226
rect 550118 514046 550174 514102
rect 550242 514046 550298 514102
rect 550118 513922 550174 513978
rect 550242 513922 550298 513978
rect 12518 508294 12574 508350
rect 12642 508294 12698 508350
rect 12518 508170 12574 508226
rect 12642 508170 12698 508226
rect 12518 508046 12574 508102
rect 12642 508046 12698 508102
rect 12518 507922 12574 507978
rect 12642 507922 12698 507978
rect 43238 508294 43294 508350
rect 43362 508294 43418 508350
rect 43238 508170 43294 508226
rect 43362 508170 43418 508226
rect 43238 508046 43294 508102
rect 43362 508046 43418 508102
rect 43238 507922 43294 507978
rect 43362 507922 43418 507978
rect 73958 508294 74014 508350
rect 74082 508294 74138 508350
rect 73958 508170 74014 508226
rect 74082 508170 74138 508226
rect 73958 508046 74014 508102
rect 74082 508046 74138 508102
rect 73958 507922 74014 507978
rect 74082 507922 74138 507978
rect 104678 508294 104734 508350
rect 104802 508294 104858 508350
rect 104678 508170 104734 508226
rect 104802 508170 104858 508226
rect 104678 508046 104734 508102
rect 104802 508046 104858 508102
rect 104678 507922 104734 507978
rect 104802 507922 104858 507978
rect 135398 508294 135454 508350
rect 135522 508294 135578 508350
rect 135398 508170 135454 508226
rect 135522 508170 135578 508226
rect 135398 508046 135454 508102
rect 135522 508046 135578 508102
rect 135398 507922 135454 507978
rect 135522 507922 135578 507978
rect 166118 508294 166174 508350
rect 166242 508294 166298 508350
rect 166118 508170 166174 508226
rect 166242 508170 166298 508226
rect 166118 508046 166174 508102
rect 166242 508046 166298 508102
rect 166118 507922 166174 507978
rect 166242 507922 166298 507978
rect 196838 508294 196894 508350
rect 196962 508294 197018 508350
rect 196838 508170 196894 508226
rect 196962 508170 197018 508226
rect 196838 508046 196894 508102
rect 196962 508046 197018 508102
rect 196838 507922 196894 507978
rect 196962 507922 197018 507978
rect 227558 508294 227614 508350
rect 227682 508294 227738 508350
rect 227558 508170 227614 508226
rect 227682 508170 227738 508226
rect 227558 508046 227614 508102
rect 227682 508046 227738 508102
rect 227558 507922 227614 507978
rect 227682 507922 227738 507978
rect 258278 508294 258334 508350
rect 258402 508294 258458 508350
rect 258278 508170 258334 508226
rect 258402 508170 258458 508226
rect 258278 508046 258334 508102
rect 258402 508046 258458 508102
rect 258278 507922 258334 507978
rect 258402 507922 258458 507978
rect 288998 508294 289054 508350
rect 289122 508294 289178 508350
rect 288998 508170 289054 508226
rect 289122 508170 289178 508226
rect 288998 508046 289054 508102
rect 289122 508046 289178 508102
rect 288998 507922 289054 507978
rect 289122 507922 289178 507978
rect 319718 508294 319774 508350
rect 319842 508294 319898 508350
rect 319718 508170 319774 508226
rect 319842 508170 319898 508226
rect 319718 508046 319774 508102
rect 319842 508046 319898 508102
rect 319718 507922 319774 507978
rect 319842 507922 319898 507978
rect 350438 508294 350494 508350
rect 350562 508294 350618 508350
rect 350438 508170 350494 508226
rect 350562 508170 350618 508226
rect 350438 508046 350494 508102
rect 350562 508046 350618 508102
rect 350438 507922 350494 507978
rect 350562 507922 350618 507978
rect 381158 508294 381214 508350
rect 381282 508294 381338 508350
rect 381158 508170 381214 508226
rect 381282 508170 381338 508226
rect 381158 508046 381214 508102
rect 381282 508046 381338 508102
rect 381158 507922 381214 507978
rect 381282 507922 381338 507978
rect 411878 508294 411934 508350
rect 412002 508294 412058 508350
rect 411878 508170 411934 508226
rect 412002 508170 412058 508226
rect 411878 508046 411934 508102
rect 412002 508046 412058 508102
rect 411878 507922 411934 507978
rect 412002 507922 412058 507978
rect 442598 508294 442654 508350
rect 442722 508294 442778 508350
rect 442598 508170 442654 508226
rect 442722 508170 442778 508226
rect 442598 508046 442654 508102
rect 442722 508046 442778 508102
rect 442598 507922 442654 507978
rect 442722 507922 442778 507978
rect 473318 508294 473374 508350
rect 473442 508294 473498 508350
rect 473318 508170 473374 508226
rect 473442 508170 473498 508226
rect 473318 508046 473374 508102
rect 473442 508046 473498 508102
rect 473318 507922 473374 507978
rect 473442 507922 473498 507978
rect 504038 508294 504094 508350
rect 504162 508294 504218 508350
rect 504038 508170 504094 508226
rect 504162 508170 504218 508226
rect 504038 508046 504094 508102
rect 504162 508046 504218 508102
rect 504038 507922 504094 507978
rect 504162 507922 504218 507978
rect 534758 508294 534814 508350
rect 534882 508294 534938 508350
rect 534758 508170 534814 508226
rect 534882 508170 534938 508226
rect 534758 508046 534814 508102
rect 534882 508046 534938 508102
rect 534758 507922 534814 507978
rect 534882 507922 534938 507978
rect 565478 508294 565534 508350
rect 565602 508294 565658 508350
rect 565478 508170 565534 508226
rect 565602 508170 565658 508226
rect 565478 508046 565534 508102
rect 565602 508046 565658 508102
rect 565478 507922 565534 507978
rect 565602 507922 565658 507978
rect 27878 496294 27934 496350
rect 28002 496294 28058 496350
rect 27878 496170 27934 496226
rect 28002 496170 28058 496226
rect 27878 496046 27934 496102
rect 28002 496046 28058 496102
rect 27878 495922 27934 495978
rect 28002 495922 28058 495978
rect 58598 496294 58654 496350
rect 58722 496294 58778 496350
rect 58598 496170 58654 496226
rect 58722 496170 58778 496226
rect 58598 496046 58654 496102
rect 58722 496046 58778 496102
rect 58598 495922 58654 495978
rect 58722 495922 58778 495978
rect 89318 496294 89374 496350
rect 89442 496294 89498 496350
rect 89318 496170 89374 496226
rect 89442 496170 89498 496226
rect 89318 496046 89374 496102
rect 89442 496046 89498 496102
rect 89318 495922 89374 495978
rect 89442 495922 89498 495978
rect 120038 496294 120094 496350
rect 120162 496294 120218 496350
rect 120038 496170 120094 496226
rect 120162 496170 120218 496226
rect 120038 496046 120094 496102
rect 120162 496046 120218 496102
rect 120038 495922 120094 495978
rect 120162 495922 120218 495978
rect 150758 496294 150814 496350
rect 150882 496294 150938 496350
rect 150758 496170 150814 496226
rect 150882 496170 150938 496226
rect 150758 496046 150814 496102
rect 150882 496046 150938 496102
rect 150758 495922 150814 495978
rect 150882 495922 150938 495978
rect 181478 496294 181534 496350
rect 181602 496294 181658 496350
rect 181478 496170 181534 496226
rect 181602 496170 181658 496226
rect 181478 496046 181534 496102
rect 181602 496046 181658 496102
rect 181478 495922 181534 495978
rect 181602 495922 181658 495978
rect 212198 496294 212254 496350
rect 212322 496294 212378 496350
rect 212198 496170 212254 496226
rect 212322 496170 212378 496226
rect 212198 496046 212254 496102
rect 212322 496046 212378 496102
rect 212198 495922 212254 495978
rect 212322 495922 212378 495978
rect 242918 496294 242974 496350
rect 243042 496294 243098 496350
rect 242918 496170 242974 496226
rect 243042 496170 243098 496226
rect 242918 496046 242974 496102
rect 243042 496046 243098 496102
rect 242918 495922 242974 495978
rect 243042 495922 243098 495978
rect 273638 496294 273694 496350
rect 273762 496294 273818 496350
rect 273638 496170 273694 496226
rect 273762 496170 273818 496226
rect 273638 496046 273694 496102
rect 273762 496046 273818 496102
rect 273638 495922 273694 495978
rect 273762 495922 273818 495978
rect 304358 496294 304414 496350
rect 304482 496294 304538 496350
rect 304358 496170 304414 496226
rect 304482 496170 304538 496226
rect 304358 496046 304414 496102
rect 304482 496046 304538 496102
rect 304358 495922 304414 495978
rect 304482 495922 304538 495978
rect 335078 496294 335134 496350
rect 335202 496294 335258 496350
rect 335078 496170 335134 496226
rect 335202 496170 335258 496226
rect 335078 496046 335134 496102
rect 335202 496046 335258 496102
rect 335078 495922 335134 495978
rect 335202 495922 335258 495978
rect 365798 496294 365854 496350
rect 365922 496294 365978 496350
rect 365798 496170 365854 496226
rect 365922 496170 365978 496226
rect 365798 496046 365854 496102
rect 365922 496046 365978 496102
rect 365798 495922 365854 495978
rect 365922 495922 365978 495978
rect 396518 496294 396574 496350
rect 396642 496294 396698 496350
rect 396518 496170 396574 496226
rect 396642 496170 396698 496226
rect 396518 496046 396574 496102
rect 396642 496046 396698 496102
rect 396518 495922 396574 495978
rect 396642 495922 396698 495978
rect 427238 496294 427294 496350
rect 427362 496294 427418 496350
rect 427238 496170 427294 496226
rect 427362 496170 427418 496226
rect 427238 496046 427294 496102
rect 427362 496046 427418 496102
rect 427238 495922 427294 495978
rect 427362 495922 427418 495978
rect 457958 496294 458014 496350
rect 458082 496294 458138 496350
rect 457958 496170 458014 496226
rect 458082 496170 458138 496226
rect 457958 496046 458014 496102
rect 458082 496046 458138 496102
rect 457958 495922 458014 495978
rect 458082 495922 458138 495978
rect 488678 496294 488734 496350
rect 488802 496294 488858 496350
rect 488678 496170 488734 496226
rect 488802 496170 488858 496226
rect 488678 496046 488734 496102
rect 488802 496046 488858 496102
rect 488678 495922 488734 495978
rect 488802 495922 488858 495978
rect 519398 496294 519454 496350
rect 519522 496294 519578 496350
rect 519398 496170 519454 496226
rect 519522 496170 519578 496226
rect 519398 496046 519454 496102
rect 519522 496046 519578 496102
rect 519398 495922 519454 495978
rect 519522 495922 519578 495978
rect 550118 496294 550174 496350
rect 550242 496294 550298 496350
rect 550118 496170 550174 496226
rect 550242 496170 550298 496226
rect 550118 496046 550174 496102
rect 550242 496046 550298 496102
rect 550118 495922 550174 495978
rect 550242 495922 550298 495978
rect 5514 490294 5570 490350
rect 5638 490294 5694 490350
rect 5762 490294 5818 490350
rect 5886 490294 5942 490350
rect 5514 490170 5570 490226
rect 5638 490170 5694 490226
rect 5762 490170 5818 490226
rect 5886 490170 5942 490226
rect 5514 490046 5570 490102
rect 5638 490046 5694 490102
rect 5762 490046 5818 490102
rect 5886 490046 5942 490102
rect 5514 489922 5570 489978
rect 5638 489922 5694 489978
rect 5762 489922 5818 489978
rect 5886 489922 5942 489978
rect -860 472294 -804 472350
rect -736 472294 -680 472350
rect -612 472294 -556 472350
rect -488 472294 -432 472350
rect -860 472170 -804 472226
rect -736 472170 -680 472226
rect -612 472170 -556 472226
rect -488 472170 -432 472226
rect -860 472046 -804 472102
rect -736 472046 -680 472102
rect -612 472046 -556 472102
rect -488 472046 -432 472102
rect -860 471922 -804 471978
rect -736 471922 -680 471978
rect -612 471922 -556 471978
rect -488 471922 -432 471978
rect 12518 490294 12574 490350
rect 12642 490294 12698 490350
rect 12518 490170 12574 490226
rect 12642 490170 12698 490226
rect 12518 490046 12574 490102
rect 12642 490046 12698 490102
rect 12518 489922 12574 489978
rect 12642 489922 12698 489978
rect 43238 490294 43294 490350
rect 43362 490294 43418 490350
rect 43238 490170 43294 490226
rect 43362 490170 43418 490226
rect 43238 490046 43294 490102
rect 43362 490046 43418 490102
rect 43238 489922 43294 489978
rect 43362 489922 43418 489978
rect 73958 490294 74014 490350
rect 74082 490294 74138 490350
rect 73958 490170 74014 490226
rect 74082 490170 74138 490226
rect 73958 490046 74014 490102
rect 74082 490046 74138 490102
rect 73958 489922 74014 489978
rect 74082 489922 74138 489978
rect 104678 490294 104734 490350
rect 104802 490294 104858 490350
rect 104678 490170 104734 490226
rect 104802 490170 104858 490226
rect 104678 490046 104734 490102
rect 104802 490046 104858 490102
rect 104678 489922 104734 489978
rect 104802 489922 104858 489978
rect 135398 490294 135454 490350
rect 135522 490294 135578 490350
rect 135398 490170 135454 490226
rect 135522 490170 135578 490226
rect 135398 490046 135454 490102
rect 135522 490046 135578 490102
rect 135398 489922 135454 489978
rect 135522 489922 135578 489978
rect 166118 490294 166174 490350
rect 166242 490294 166298 490350
rect 166118 490170 166174 490226
rect 166242 490170 166298 490226
rect 166118 490046 166174 490102
rect 166242 490046 166298 490102
rect 166118 489922 166174 489978
rect 166242 489922 166298 489978
rect 196838 490294 196894 490350
rect 196962 490294 197018 490350
rect 196838 490170 196894 490226
rect 196962 490170 197018 490226
rect 196838 490046 196894 490102
rect 196962 490046 197018 490102
rect 196838 489922 196894 489978
rect 196962 489922 197018 489978
rect 227558 490294 227614 490350
rect 227682 490294 227738 490350
rect 227558 490170 227614 490226
rect 227682 490170 227738 490226
rect 227558 490046 227614 490102
rect 227682 490046 227738 490102
rect 227558 489922 227614 489978
rect 227682 489922 227738 489978
rect 258278 490294 258334 490350
rect 258402 490294 258458 490350
rect 258278 490170 258334 490226
rect 258402 490170 258458 490226
rect 258278 490046 258334 490102
rect 258402 490046 258458 490102
rect 258278 489922 258334 489978
rect 258402 489922 258458 489978
rect 288998 490294 289054 490350
rect 289122 490294 289178 490350
rect 288998 490170 289054 490226
rect 289122 490170 289178 490226
rect 288998 490046 289054 490102
rect 289122 490046 289178 490102
rect 288998 489922 289054 489978
rect 289122 489922 289178 489978
rect 319718 490294 319774 490350
rect 319842 490294 319898 490350
rect 319718 490170 319774 490226
rect 319842 490170 319898 490226
rect 319718 490046 319774 490102
rect 319842 490046 319898 490102
rect 319718 489922 319774 489978
rect 319842 489922 319898 489978
rect 350438 490294 350494 490350
rect 350562 490294 350618 490350
rect 350438 490170 350494 490226
rect 350562 490170 350618 490226
rect 350438 490046 350494 490102
rect 350562 490046 350618 490102
rect 350438 489922 350494 489978
rect 350562 489922 350618 489978
rect 381158 490294 381214 490350
rect 381282 490294 381338 490350
rect 381158 490170 381214 490226
rect 381282 490170 381338 490226
rect 381158 490046 381214 490102
rect 381282 490046 381338 490102
rect 381158 489922 381214 489978
rect 381282 489922 381338 489978
rect 411878 490294 411934 490350
rect 412002 490294 412058 490350
rect 411878 490170 411934 490226
rect 412002 490170 412058 490226
rect 411878 490046 411934 490102
rect 412002 490046 412058 490102
rect 411878 489922 411934 489978
rect 412002 489922 412058 489978
rect 442598 490294 442654 490350
rect 442722 490294 442778 490350
rect 442598 490170 442654 490226
rect 442722 490170 442778 490226
rect 442598 490046 442654 490102
rect 442722 490046 442778 490102
rect 442598 489922 442654 489978
rect 442722 489922 442778 489978
rect 473318 490294 473374 490350
rect 473442 490294 473498 490350
rect 473318 490170 473374 490226
rect 473442 490170 473498 490226
rect 473318 490046 473374 490102
rect 473442 490046 473498 490102
rect 473318 489922 473374 489978
rect 473442 489922 473498 489978
rect 504038 490294 504094 490350
rect 504162 490294 504218 490350
rect 504038 490170 504094 490226
rect 504162 490170 504218 490226
rect 504038 490046 504094 490102
rect 504162 490046 504218 490102
rect 504038 489922 504094 489978
rect 504162 489922 504218 489978
rect 534758 490294 534814 490350
rect 534882 490294 534938 490350
rect 534758 490170 534814 490226
rect 534882 490170 534938 490226
rect 534758 490046 534814 490102
rect 534882 490046 534938 490102
rect 534758 489922 534814 489978
rect 534882 489922 534938 489978
rect 565478 490294 565534 490350
rect 565602 490294 565658 490350
rect 589194 508294 589250 508350
rect 589318 508294 589374 508350
rect 589442 508294 589498 508350
rect 589566 508294 589622 508350
rect 589194 508170 589250 508226
rect 589318 508170 589374 508226
rect 589442 508170 589498 508226
rect 589566 508170 589622 508226
rect 589194 508046 589250 508102
rect 589318 508046 589374 508102
rect 589442 508046 589498 508102
rect 589566 508046 589622 508102
rect 589194 507922 589250 507978
rect 589318 507922 589374 507978
rect 589442 507922 589498 507978
rect 589566 507922 589622 507978
rect 592914 532294 592970 532350
rect 593038 532294 593094 532350
rect 593162 532294 593218 532350
rect 593286 532294 593342 532350
rect 592914 532170 592970 532226
rect 593038 532170 593094 532226
rect 593162 532170 593218 532226
rect 593286 532170 593342 532226
rect 592914 532046 592970 532102
rect 593038 532046 593094 532102
rect 593162 532046 593218 532102
rect 593286 532046 593342 532102
rect 592914 531922 592970 531978
rect 593038 531922 593094 531978
rect 593162 531922 593218 531978
rect 593286 531922 593342 531978
rect 592914 514294 592970 514350
rect 593038 514294 593094 514350
rect 593162 514294 593218 514350
rect 593286 514294 593342 514350
rect 592914 514170 592970 514226
rect 593038 514170 593094 514226
rect 593162 514170 593218 514226
rect 593286 514170 593342 514226
rect 592914 514046 592970 514102
rect 593038 514046 593094 514102
rect 593162 514046 593218 514102
rect 593286 514046 593342 514102
rect 592914 513922 592970 513978
rect 593038 513922 593094 513978
rect 593162 513922 593218 513978
rect 593286 513922 593342 513978
rect 592914 496294 592970 496350
rect 593038 496294 593094 496350
rect 593162 496294 593218 496350
rect 593286 496294 593342 496350
rect 592914 496170 592970 496226
rect 593038 496170 593094 496226
rect 593162 496170 593218 496226
rect 593286 496170 593342 496226
rect 589194 490294 589250 490350
rect 589318 490294 589374 490350
rect 589442 490294 589498 490350
rect 589566 490294 589622 490350
rect 565478 490170 565534 490226
rect 565602 490170 565658 490226
rect 565478 490046 565534 490102
rect 565602 490046 565658 490102
rect 565478 489922 565534 489978
rect 565602 489922 565658 489978
rect 589194 490170 589250 490226
rect 589318 490170 589374 490226
rect 589442 490170 589498 490226
rect 589566 490170 589622 490226
rect 589194 490046 589250 490102
rect 589318 490046 589374 490102
rect 589442 490046 589498 490102
rect 589566 490046 589622 490102
rect 589194 489922 589250 489978
rect 589318 489922 589374 489978
rect 589442 489922 589498 489978
rect 589566 489922 589622 489978
rect 27878 478294 27934 478350
rect 28002 478294 28058 478350
rect 27878 478170 27934 478226
rect 28002 478170 28058 478226
rect 27878 478046 27934 478102
rect 28002 478046 28058 478102
rect 27878 477922 27934 477978
rect 28002 477922 28058 477978
rect 58598 478294 58654 478350
rect 58722 478294 58778 478350
rect 58598 478170 58654 478226
rect 58722 478170 58778 478226
rect 58598 478046 58654 478102
rect 58722 478046 58778 478102
rect 58598 477922 58654 477978
rect 58722 477922 58778 477978
rect 89318 478294 89374 478350
rect 89442 478294 89498 478350
rect 89318 478170 89374 478226
rect 89442 478170 89498 478226
rect 89318 478046 89374 478102
rect 89442 478046 89498 478102
rect 89318 477922 89374 477978
rect 89442 477922 89498 477978
rect 120038 478294 120094 478350
rect 120162 478294 120218 478350
rect 120038 478170 120094 478226
rect 120162 478170 120218 478226
rect 120038 478046 120094 478102
rect 120162 478046 120218 478102
rect 120038 477922 120094 477978
rect 120162 477922 120218 477978
rect 150758 478294 150814 478350
rect 150882 478294 150938 478350
rect 150758 478170 150814 478226
rect 150882 478170 150938 478226
rect 150758 478046 150814 478102
rect 150882 478046 150938 478102
rect 150758 477922 150814 477978
rect 150882 477922 150938 477978
rect 181478 478294 181534 478350
rect 181602 478294 181658 478350
rect 181478 478170 181534 478226
rect 181602 478170 181658 478226
rect 181478 478046 181534 478102
rect 181602 478046 181658 478102
rect 181478 477922 181534 477978
rect 181602 477922 181658 477978
rect 212198 478294 212254 478350
rect 212322 478294 212378 478350
rect 212198 478170 212254 478226
rect 212322 478170 212378 478226
rect 212198 478046 212254 478102
rect 212322 478046 212378 478102
rect 212198 477922 212254 477978
rect 212322 477922 212378 477978
rect 242918 478294 242974 478350
rect 243042 478294 243098 478350
rect 242918 478170 242974 478226
rect 243042 478170 243098 478226
rect 242918 478046 242974 478102
rect 243042 478046 243098 478102
rect 242918 477922 242974 477978
rect 243042 477922 243098 477978
rect 273638 478294 273694 478350
rect 273762 478294 273818 478350
rect 273638 478170 273694 478226
rect 273762 478170 273818 478226
rect 273638 478046 273694 478102
rect 273762 478046 273818 478102
rect 273638 477922 273694 477978
rect 273762 477922 273818 477978
rect 304358 478294 304414 478350
rect 304482 478294 304538 478350
rect 304358 478170 304414 478226
rect 304482 478170 304538 478226
rect 304358 478046 304414 478102
rect 304482 478046 304538 478102
rect 304358 477922 304414 477978
rect 304482 477922 304538 477978
rect 335078 478294 335134 478350
rect 335202 478294 335258 478350
rect 335078 478170 335134 478226
rect 335202 478170 335258 478226
rect 335078 478046 335134 478102
rect 335202 478046 335258 478102
rect 335078 477922 335134 477978
rect 335202 477922 335258 477978
rect 365798 478294 365854 478350
rect 365922 478294 365978 478350
rect 365798 478170 365854 478226
rect 365922 478170 365978 478226
rect 365798 478046 365854 478102
rect 365922 478046 365978 478102
rect 365798 477922 365854 477978
rect 365922 477922 365978 477978
rect 396518 478294 396574 478350
rect 396642 478294 396698 478350
rect 396518 478170 396574 478226
rect 396642 478170 396698 478226
rect 396518 478046 396574 478102
rect 396642 478046 396698 478102
rect 396518 477922 396574 477978
rect 396642 477922 396698 477978
rect 427238 478294 427294 478350
rect 427362 478294 427418 478350
rect 427238 478170 427294 478226
rect 427362 478170 427418 478226
rect 427238 478046 427294 478102
rect 427362 478046 427418 478102
rect 427238 477922 427294 477978
rect 427362 477922 427418 477978
rect 457958 478294 458014 478350
rect 458082 478294 458138 478350
rect 457958 478170 458014 478226
rect 458082 478170 458138 478226
rect 457958 478046 458014 478102
rect 458082 478046 458138 478102
rect 457958 477922 458014 477978
rect 458082 477922 458138 477978
rect 488678 478294 488734 478350
rect 488802 478294 488858 478350
rect 488678 478170 488734 478226
rect 488802 478170 488858 478226
rect 488678 478046 488734 478102
rect 488802 478046 488858 478102
rect 488678 477922 488734 477978
rect 488802 477922 488858 477978
rect 519398 478294 519454 478350
rect 519522 478294 519578 478350
rect 519398 478170 519454 478226
rect 519522 478170 519578 478226
rect 519398 478046 519454 478102
rect 519522 478046 519578 478102
rect 519398 477922 519454 477978
rect 519522 477922 519578 477978
rect 550118 478294 550174 478350
rect 550242 478294 550298 478350
rect 550118 478170 550174 478226
rect 550242 478170 550298 478226
rect 550118 478046 550174 478102
rect 550242 478046 550298 478102
rect 550118 477922 550174 477978
rect 550242 477922 550298 477978
rect 5514 472294 5570 472350
rect 5638 472294 5694 472350
rect 5762 472294 5818 472350
rect 5886 472294 5942 472350
rect 5514 472170 5570 472226
rect 5638 472170 5694 472226
rect 5762 472170 5818 472226
rect 5886 472170 5942 472226
rect 5514 472046 5570 472102
rect 5638 472046 5694 472102
rect 5762 472046 5818 472102
rect 5886 472046 5942 472102
rect 5514 471922 5570 471978
rect 5638 471922 5694 471978
rect 5762 471922 5818 471978
rect 5886 471922 5942 471978
rect -860 454294 -804 454350
rect -736 454294 -680 454350
rect -612 454294 -556 454350
rect -488 454294 -432 454350
rect -860 454170 -804 454226
rect -736 454170 -680 454226
rect -612 454170 -556 454226
rect -488 454170 -432 454226
rect -860 454046 -804 454102
rect -736 454046 -680 454102
rect -612 454046 -556 454102
rect -488 454046 -432 454102
rect -860 453922 -804 453978
rect -736 453922 -680 453978
rect -612 453922 -556 453978
rect -488 453922 -432 453978
rect 5514 454294 5570 454350
rect 5638 454294 5694 454350
rect 5762 454294 5818 454350
rect 5886 454294 5942 454350
rect 5514 454170 5570 454226
rect 5638 454170 5694 454226
rect 5762 454170 5818 454226
rect 5886 454170 5942 454226
rect 5514 454046 5570 454102
rect 5638 454046 5694 454102
rect 5762 454046 5818 454102
rect 5886 454046 5942 454102
rect 5514 453922 5570 453978
rect 5638 453922 5694 453978
rect 5762 453922 5818 453978
rect 5886 453922 5942 453978
rect -860 436294 -804 436350
rect -736 436294 -680 436350
rect -612 436294 -556 436350
rect -488 436294 -432 436350
rect -860 436170 -804 436226
rect -736 436170 -680 436226
rect -612 436170 -556 436226
rect -488 436170 -432 436226
rect -860 436046 -804 436102
rect -736 436046 -680 436102
rect -612 436046 -556 436102
rect -488 436046 -432 436102
rect -860 435922 -804 435978
rect -736 435922 -680 435978
rect -612 435922 -556 435978
rect -488 435922 -432 435978
rect 12518 472294 12574 472350
rect 12642 472294 12698 472350
rect 12518 472170 12574 472226
rect 12642 472170 12698 472226
rect 12518 472046 12574 472102
rect 12642 472046 12698 472102
rect 12518 471922 12574 471978
rect 12642 471922 12698 471978
rect 43238 472294 43294 472350
rect 43362 472294 43418 472350
rect 43238 472170 43294 472226
rect 43362 472170 43418 472226
rect 43238 472046 43294 472102
rect 43362 472046 43418 472102
rect 43238 471922 43294 471978
rect 43362 471922 43418 471978
rect 73958 472294 74014 472350
rect 74082 472294 74138 472350
rect 73958 472170 74014 472226
rect 74082 472170 74138 472226
rect 73958 472046 74014 472102
rect 74082 472046 74138 472102
rect 73958 471922 74014 471978
rect 74082 471922 74138 471978
rect 104678 472294 104734 472350
rect 104802 472294 104858 472350
rect 104678 472170 104734 472226
rect 104802 472170 104858 472226
rect 104678 472046 104734 472102
rect 104802 472046 104858 472102
rect 104678 471922 104734 471978
rect 104802 471922 104858 471978
rect 135398 472294 135454 472350
rect 135522 472294 135578 472350
rect 135398 472170 135454 472226
rect 135522 472170 135578 472226
rect 135398 472046 135454 472102
rect 135522 472046 135578 472102
rect 135398 471922 135454 471978
rect 135522 471922 135578 471978
rect 166118 472294 166174 472350
rect 166242 472294 166298 472350
rect 166118 472170 166174 472226
rect 166242 472170 166298 472226
rect 166118 472046 166174 472102
rect 166242 472046 166298 472102
rect 166118 471922 166174 471978
rect 166242 471922 166298 471978
rect 196838 472294 196894 472350
rect 196962 472294 197018 472350
rect 196838 472170 196894 472226
rect 196962 472170 197018 472226
rect 196838 472046 196894 472102
rect 196962 472046 197018 472102
rect 196838 471922 196894 471978
rect 196962 471922 197018 471978
rect 227558 472294 227614 472350
rect 227682 472294 227738 472350
rect 227558 472170 227614 472226
rect 227682 472170 227738 472226
rect 227558 472046 227614 472102
rect 227682 472046 227738 472102
rect 227558 471922 227614 471978
rect 227682 471922 227738 471978
rect 258278 472294 258334 472350
rect 258402 472294 258458 472350
rect 258278 472170 258334 472226
rect 258402 472170 258458 472226
rect 258278 472046 258334 472102
rect 258402 472046 258458 472102
rect 258278 471922 258334 471978
rect 258402 471922 258458 471978
rect 288998 472294 289054 472350
rect 289122 472294 289178 472350
rect 288998 472170 289054 472226
rect 289122 472170 289178 472226
rect 288998 472046 289054 472102
rect 289122 472046 289178 472102
rect 288998 471922 289054 471978
rect 289122 471922 289178 471978
rect 319718 472294 319774 472350
rect 319842 472294 319898 472350
rect 319718 472170 319774 472226
rect 319842 472170 319898 472226
rect 319718 472046 319774 472102
rect 319842 472046 319898 472102
rect 319718 471922 319774 471978
rect 319842 471922 319898 471978
rect 350438 472294 350494 472350
rect 350562 472294 350618 472350
rect 350438 472170 350494 472226
rect 350562 472170 350618 472226
rect 350438 472046 350494 472102
rect 350562 472046 350618 472102
rect 350438 471922 350494 471978
rect 350562 471922 350618 471978
rect 381158 472294 381214 472350
rect 381282 472294 381338 472350
rect 381158 472170 381214 472226
rect 381282 472170 381338 472226
rect 381158 472046 381214 472102
rect 381282 472046 381338 472102
rect 381158 471922 381214 471978
rect 381282 471922 381338 471978
rect 411878 472294 411934 472350
rect 412002 472294 412058 472350
rect 411878 472170 411934 472226
rect 412002 472170 412058 472226
rect 411878 472046 411934 472102
rect 412002 472046 412058 472102
rect 411878 471922 411934 471978
rect 412002 471922 412058 471978
rect 442598 472294 442654 472350
rect 442722 472294 442778 472350
rect 442598 472170 442654 472226
rect 442722 472170 442778 472226
rect 442598 472046 442654 472102
rect 442722 472046 442778 472102
rect 442598 471922 442654 471978
rect 442722 471922 442778 471978
rect 473318 472294 473374 472350
rect 473442 472294 473498 472350
rect 473318 472170 473374 472226
rect 473442 472170 473498 472226
rect 473318 472046 473374 472102
rect 473442 472046 473498 472102
rect 473318 471922 473374 471978
rect 473442 471922 473498 471978
rect 504038 472294 504094 472350
rect 504162 472294 504218 472350
rect 504038 472170 504094 472226
rect 504162 472170 504218 472226
rect 504038 472046 504094 472102
rect 504162 472046 504218 472102
rect 504038 471922 504094 471978
rect 504162 471922 504218 471978
rect 534758 472294 534814 472350
rect 534882 472294 534938 472350
rect 534758 472170 534814 472226
rect 534882 472170 534938 472226
rect 534758 472046 534814 472102
rect 534882 472046 534938 472102
rect 534758 471922 534814 471978
rect 534882 471922 534938 471978
rect 565478 472294 565534 472350
rect 565602 472294 565658 472350
rect 565478 472170 565534 472226
rect 565602 472170 565658 472226
rect 565478 472046 565534 472102
rect 565602 472046 565658 472102
rect 565478 471922 565534 471978
rect 565602 471922 565658 471978
rect 592914 496046 592970 496102
rect 593038 496046 593094 496102
rect 593162 496046 593218 496102
rect 593286 496046 593342 496102
rect 592914 495922 592970 495978
rect 593038 495922 593094 495978
rect 593162 495922 593218 495978
rect 593286 495922 593342 495978
rect 589194 472294 589250 472350
rect 589318 472294 589374 472350
rect 589442 472294 589498 472350
rect 589566 472294 589622 472350
rect 589194 472170 589250 472226
rect 589318 472170 589374 472226
rect 589442 472170 589498 472226
rect 589566 472170 589622 472226
rect 589194 472046 589250 472102
rect 589318 472046 589374 472102
rect 589442 472046 589498 472102
rect 589566 472046 589622 472102
rect 589194 471922 589250 471978
rect 589318 471922 589374 471978
rect 589442 471922 589498 471978
rect 589566 471922 589622 471978
rect 27878 460294 27934 460350
rect 28002 460294 28058 460350
rect 27878 460170 27934 460226
rect 28002 460170 28058 460226
rect 27878 460046 27934 460102
rect 28002 460046 28058 460102
rect 27878 459922 27934 459978
rect 28002 459922 28058 459978
rect 58598 460294 58654 460350
rect 58722 460294 58778 460350
rect 58598 460170 58654 460226
rect 58722 460170 58778 460226
rect 58598 460046 58654 460102
rect 58722 460046 58778 460102
rect 58598 459922 58654 459978
rect 58722 459922 58778 459978
rect 89318 460294 89374 460350
rect 89442 460294 89498 460350
rect 89318 460170 89374 460226
rect 89442 460170 89498 460226
rect 89318 460046 89374 460102
rect 89442 460046 89498 460102
rect 89318 459922 89374 459978
rect 89442 459922 89498 459978
rect 120038 460294 120094 460350
rect 120162 460294 120218 460350
rect 120038 460170 120094 460226
rect 120162 460170 120218 460226
rect 120038 460046 120094 460102
rect 120162 460046 120218 460102
rect 120038 459922 120094 459978
rect 120162 459922 120218 459978
rect 150758 460294 150814 460350
rect 150882 460294 150938 460350
rect 150758 460170 150814 460226
rect 150882 460170 150938 460226
rect 150758 460046 150814 460102
rect 150882 460046 150938 460102
rect 150758 459922 150814 459978
rect 150882 459922 150938 459978
rect 181478 460294 181534 460350
rect 181602 460294 181658 460350
rect 181478 460170 181534 460226
rect 181602 460170 181658 460226
rect 181478 460046 181534 460102
rect 181602 460046 181658 460102
rect 181478 459922 181534 459978
rect 181602 459922 181658 459978
rect 212198 460294 212254 460350
rect 212322 460294 212378 460350
rect 212198 460170 212254 460226
rect 212322 460170 212378 460226
rect 212198 460046 212254 460102
rect 212322 460046 212378 460102
rect 212198 459922 212254 459978
rect 212322 459922 212378 459978
rect 242918 460294 242974 460350
rect 243042 460294 243098 460350
rect 242918 460170 242974 460226
rect 243042 460170 243098 460226
rect 242918 460046 242974 460102
rect 243042 460046 243098 460102
rect 242918 459922 242974 459978
rect 243042 459922 243098 459978
rect 273638 460294 273694 460350
rect 273762 460294 273818 460350
rect 273638 460170 273694 460226
rect 273762 460170 273818 460226
rect 273638 460046 273694 460102
rect 273762 460046 273818 460102
rect 273638 459922 273694 459978
rect 273762 459922 273818 459978
rect 304358 460294 304414 460350
rect 304482 460294 304538 460350
rect 304358 460170 304414 460226
rect 304482 460170 304538 460226
rect 304358 460046 304414 460102
rect 304482 460046 304538 460102
rect 304358 459922 304414 459978
rect 304482 459922 304538 459978
rect 335078 460294 335134 460350
rect 335202 460294 335258 460350
rect 335078 460170 335134 460226
rect 335202 460170 335258 460226
rect 335078 460046 335134 460102
rect 335202 460046 335258 460102
rect 335078 459922 335134 459978
rect 335202 459922 335258 459978
rect 365798 460294 365854 460350
rect 365922 460294 365978 460350
rect 365798 460170 365854 460226
rect 365922 460170 365978 460226
rect 365798 460046 365854 460102
rect 365922 460046 365978 460102
rect 365798 459922 365854 459978
rect 365922 459922 365978 459978
rect 396518 460294 396574 460350
rect 396642 460294 396698 460350
rect 396518 460170 396574 460226
rect 396642 460170 396698 460226
rect 396518 460046 396574 460102
rect 396642 460046 396698 460102
rect 396518 459922 396574 459978
rect 396642 459922 396698 459978
rect 427238 460294 427294 460350
rect 427362 460294 427418 460350
rect 427238 460170 427294 460226
rect 427362 460170 427418 460226
rect 427238 460046 427294 460102
rect 427362 460046 427418 460102
rect 427238 459922 427294 459978
rect 427362 459922 427418 459978
rect 457958 460294 458014 460350
rect 458082 460294 458138 460350
rect 457958 460170 458014 460226
rect 458082 460170 458138 460226
rect 457958 460046 458014 460102
rect 458082 460046 458138 460102
rect 457958 459922 458014 459978
rect 458082 459922 458138 459978
rect 488678 460294 488734 460350
rect 488802 460294 488858 460350
rect 488678 460170 488734 460226
rect 488802 460170 488858 460226
rect 488678 460046 488734 460102
rect 488802 460046 488858 460102
rect 488678 459922 488734 459978
rect 488802 459922 488858 459978
rect 519398 460294 519454 460350
rect 519522 460294 519578 460350
rect 519398 460170 519454 460226
rect 519522 460170 519578 460226
rect 519398 460046 519454 460102
rect 519522 460046 519578 460102
rect 519398 459922 519454 459978
rect 519522 459922 519578 459978
rect 550118 460294 550174 460350
rect 550242 460294 550298 460350
rect 550118 460170 550174 460226
rect 550242 460170 550298 460226
rect 550118 460046 550174 460102
rect 550242 460046 550298 460102
rect 550118 459922 550174 459978
rect 550242 459922 550298 459978
rect 12518 454294 12574 454350
rect 12642 454294 12698 454350
rect 12518 454170 12574 454226
rect 12642 454170 12698 454226
rect 12518 454046 12574 454102
rect 12642 454046 12698 454102
rect 12518 453922 12574 453978
rect 12642 453922 12698 453978
rect 43238 454294 43294 454350
rect 43362 454294 43418 454350
rect 43238 454170 43294 454226
rect 43362 454170 43418 454226
rect 43238 454046 43294 454102
rect 43362 454046 43418 454102
rect 43238 453922 43294 453978
rect 43362 453922 43418 453978
rect 73958 454294 74014 454350
rect 74082 454294 74138 454350
rect 73958 454170 74014 454226
rect 74082 454170 74138 454226
rect 73958 454046 74014 454102
rect 74082 454046 74138 454102
rect 73958 453922 74014 453978
rect 74082 453922 74138 453978
rect 104678 454294 104734 454350
rect 104802 454294 104858 454350
rect 104678 454170 104734 454226
rect 104802 454170 104858 454226
rect 104678 454046 104734 454102
rect 104802 454046 104858 454102
rect 104678 453922 104734 453978
rect 104802 453922 104858 453978
rect 135398 454294 135454 454350
rect 135522 454294 135578 454350
rect 135398 454170 135454 454226
rect 135522 454170 135578 454226
rect 135398 454046 135454 454102
rect 135522 454046 135578 454102
rect 135398 453922 135454 453978
rect 135522 453922 135578 453978
rect 166118 454294 166174 454350
rect 166242 454294 166298 454350
rect 166118 454170 166174 454226
rect 166242 454170 166298 454226
rect 166118 454046 166174 454102
rect 166242 454046 166298 454102
rect 166118 453922 166174 453978
rect 166242 453922 166298 453978
rect 196838 454294 196894 454350
rect 196962 454294 197018 454350
rect 196838 454170 196894 454226
rect 196962 454170 197018 454226
rect 196838 454046 196894 454102
rect 196962 454046 197018 454102
rect 196838 453922 196894 453978
rect 196962 453922 197018 453978
rect 227558 454294 227614 454350
rect 227682 454294 227738 454350
rect 227558 454170 227614 454226
rect 227682 454170 227738 454226
rect 227558 454046 227614 454102
rect 227682 454046 227738 454102
rect 227558 453922 227614 453978
rect 227682 453922 227738 453978
rect 258278 454294 258334 454350
rect 258402 454294 258458 454350
rect 258278 454170 258334 454226
rect 258402 454170 258458 454226
rect 258278 454046 258334 454102
rect 258402 454046 258458 454102
rect 258278 453922 258334 453978
rect 258402 453922 258458 453978
rect 288998 454294 289054 454350
rect 289122 454294 289178 454350
rect 288998 454170 289054 454226
rect 289122 454170 289178 454226
rect 288998 454046 289054 454102
rect 289122 454046 289178 454102
rect 288998 453922 289054 453978
rect 289122 453922 289178 453978
rect 319718 454294 319774 454350
rect 319842 454294 319898 454350
rect 319718 454170 319774 454226
rect 319842 454170 319898 454226
rect 319718 454046 319774 454102
rect 319842 454046 319898 454102
rect 319718 453922 319774 453978
rect 319842 453922 319898 453978
rect 350438 454294 350494 454350
rect 350562 454294 350618 454350
rect 350438 454170 350494 454226
rect 350562 454170 350618 454226
rect 350438 454046 350494 454102
rect 350562 454046 350618 454102
rect 350438 453922 350494 453978
rect 350562 453922 350618 453978
rect 381158 454294 381214 454350
rect 381282 454294 381338 454350
rect 381158 454170 381214 454226
rect 381282 454170 381338 454226
rect 381158 454046 381214 454102
rect 381282 454046 381338 454102
rect 381158 453922 381214 453978
rect 381282 453922 381338 453978
rect 411878 454294 411934 454350
rect 412002 454294 412058 454350
rect 411878 454170 411934 454226
rect 412002 454170 412058 454226
rect 411878 454046 411934 454102
rect 412002 454046 412058 454102
rect 411878 453922 411934 453978
rect 412002 453922 412058 453978
rect 442598 454294 442654 454350
rect 442722 454294 442778 454350
rect 442598 454170 442654 454226
rect 442722 454170 442778 454226
rect 442598 454046 442654 454102
rect 442722 454046 442778 454102
rect 442598 453922 442654 453978
rect 442722 453922 442778 453978
rect 473318 454294 473374 454350
rect 473442 454294 473498 454350
rect 473318 454170 473374 454226
rect 473442 454170 473498 454226
rect 473318 454046 473374 454102
rect 473442 454046 473498 454102
rect 473318 453922 473374 453978
rect 473442 453922 473498 453978
rect 504038 454294 504094 454350
rect 504162 454294 504218 454350
rect 504038 454170 504094 454226
rect 504162 454170 504218 454226
rect 504038 454046 504094 454102
rect 504162 454046 504218 454102
rect 504038 453922 504094 453978
rect 504162 453922 504218 453978
rect 534758 454294 534814 454350
rect 534882 454294 534938 454350
rect 534758 454170 534814 454226
rect 534882 454170 534938 454226
rect 534758 454046 534814 454102
rect 534882 454046 534938 454102
rect 534758 453922 534814 453978
rect 534882 453922 534938 453978
rect 565478 454294 565534 454350
rect 565602 454294 565658 454350
rect 565478 454170 565534 454226
rect 565602 454170 565658 454226
rect 565478 454046 565534 454102
rect 565602 454046 565658 454102
rect 565478 453922 565534 453978
rect 565602 453922 565658 453978
rect 27878 442294 27934 442350
rect 28002 442294 28058 442350
rect 27878 442170 27934 442226
rect 28002 442170 28058 442226
rect 27878 442046 27934 442102
rect 28002 442046 28058 442102
rect 27878 441922 27934 441978
rect 28002 441922 28058 441978
rect 58598 442294 58654 442350
rect 58722 442294 58778 442350
rect 58598 442170 58654 442226
rect 58722 442170 58778 442226
rect 58598 442046 58654 442102
rect 58722 442046 58778 442102
rect 58598 441922 58654 441978
rect 58722 441922 58778 441978
rect 89318 442294 89374 442350
rect 89442 442294 89498 442350
rect 89318 442170 89374 442226
rect 89442 442170 89498 442226
rect 89318 442046 89374 442102
rect 89442 442046 89498 442102
rect 89318 441922 89374 441978
rect 89442 441922 89498 441978
rect 120038 442294 120094 442350
rect 120162 442294 120218 442350
rect 120038 442170 120094 442226
rect 120162 442170 120218 442226
rect 120038 442046 120094 442102
rect 120162 442046 120218 442102
rect 120038 441922 120094 441978
rect 120162 441922 120218 441978
rect 150758 442294 150814 442350
rect 150882 442294 150938 442350
rect 150758 442170 150814 442226
rect 150882 442170 150938 442226
rect 150758 442046 150814 442102
rect 150882 442046 150938 442102
rect 150758 441922 150814 441978
rect 150882 441922 150938 441978
rect 181478 442294 181534 442350
rect 181602 442294 181658 442350
rect 181478 442170 181534 442226
rect 181602 442170 181658 442226
rect 181478 442046 181534 442102
rect 181602 442046 181658 442102
rect 181478 441922 181534 441978
rect 181602 441922 181658 441978
rect 212198 442294 212254 442350
rect 212322 442294 212378 442350
rect 212198 442170 212254 442226
rect 212322 442170 212378 442226
rect 212198 442046 212254 442102
rect 212322 442046 212378 442102
rect 212198 441922 212254 441978
rect 212322 441922 212378 441978
rect 242918 442294 242974 442350
rect 243042 442294 243098 442350
rect 242918 442170 242974 442226
rect 243042 442170 243098 442226
rect 242918 442046 242974 442102
rect 243042 442046 243098 442102
rect 242918 441922 242974 441978
rect 243042 441922 243098 441978
rect 273638 442294 273694 442350
rect 273762 442294 273818 442350
rect 273638 442170 273694 442226
rect 273762 442170 273818 442226
rect 273638 442046 273694 442102
rect 273762 442046 273818 442102
rect 273638 441922 273694 441978
rect 273762 441922 273818 441978
rect 304358 442294 304414 442350
rect 304482 442294 304538 442350
rect 304358 442170 304414 442226
rect 304482 442170 304538 442226
rect 304358 442046 304414 442102
rect 304482 442046 304538 442102
rect 304358 441922 304414 441978
rect 304482 441922 304538 441978
rect 335078 442294 335134 442350
rect 335202 442294 335258 442350
rect 335078 442170 335134 442226
rect 335202 442170 335258 442226
rect 335078 442046 335134 442102
rect 335202 442046 335258 442102
rect 335078 441922 335134 441978
rect 335202 441922 335258 441978
rect 365798 442294 365854 442350
rect 365922 442294 365978 442350
rect 365798 442170 365854 442226
rect 365922 442170 365978 442226
rect 365798 442046 365854 442102
rect 365922 442046 365978 442102
rect 365798 441922 365854 441978
rect 365922 441922 365978 441978
rect 396518 442294 396574 442350
rect 396642 442294 396698 442350
rect 396518 442170 396574 442226
rect 396642 442170 396698 442226
rect 396518 442046 396574 442102
rect 396642 442046 396698 442102
rect 396518 441922 396574 441978
rect 396642 441922 396698 441978
rect 427238 442294 427294 442350
rect 427362 442294 427418 442350
rect 427238 442170 427294 442226
rect 427362 442170 427418 442226
rect 427238 442046 427294 442102
rect 427362 442046 427418 442102
rect 427238 441922 427294 441978
rect 427362 441922 427418 441978
rect 457958 442294 458014 442350
rect 458082 442294 458138 442350
rect 457958 442170 458014 442226
rect 458082 442170 458138 442226
rect 457958 442046 458014 442102
rect 458082 442046 458138 442102
rect 457958 441922 458014 441978
rect 458082 441922 458138 441978
rect 488678 442294 488734 442350
rect 488802 442294 488858 442350
rect 488678 442170 488734 442226
rect 488802 442170 488858 442226
rect 488678 442046 488734 442102
rect 488802 442046 488858 442102
rect 488678 441922 488734 441978
rect 488802 441922 488858 441978
rect 519398 442294 519454 442350
rect 519522 442294 519578 442350
rect 519398 442170 519454 442226
rect 519522 442170 519578 442226
rect 519398 442046 519454 442102
rect 519522 442046 519578 442102
rect 519398 441922 519454 441978
rect 519522 441922 519578 441978
rect 550118 442294 550174 442350
rect 550242 442294 550298 442350
rect 550118 442170 550174 442226
rect 550242 442170 550298 442226
rect 550118 442046 550174 442102
rect 550242 442046 550298 442102
rect 550118 441922 550174 441978
rect 550242 441922 550298 441978
rect 592914 478294 592970 478350
rect 593038 478294 593094 478350
rect 593162 478294 593218 478350
rect 593286 478294 593342 478350
rect 592914 478170 592970 478226
rect 593038 478170 593094 478226
rect 593162 478170 593218 478226
rect 593286 478170 593342 478226
rect 592914 478046 592970 478102
rect 593038 478046 593094 478102
rect 593162 478046 593218 478102
rect 593286 478046 593342 478102
rect 592914 477922 592970 477978
rect 593038 477922 593094 477978
rect 593162 477922 593218 477978
rect 593286 477922 593342 477978
rect 589194 454294 589250 454350
rect 589318 454294 589374 454350
rect 589442 454294 589498 454350
rect 589566 454294 589622 454350
rect 589194 454170 589250 454226
rect 589318 454170 589374 454226
rect 589442 454170 589498 454226
rect 589566 454170 589622 454226
rect 589194 454046 589250 454102
rect 589318 454046 589374 454102
rect 589442 454046 589498 454102
rect 589566 454046 589622 454102
rect 589194 453922 589250 453978
rect 589318 453922 589374 453978
rect 589442 453922 589498 453978
rect 589566 453922 589622 453978
rect 5514 436294 5570 436350
rect 5638 436294 5694 436350
rect 5762 436294 5818 436350
rect 5886 436294 5942 436350
rect 5514 436170 5570 436226
rect 5638 436170 5694 436226
rect 5762 436170 5818 436226
rect 5886 436170 5942 436226
rect 5514 436046 5570 436102
rect 5638 436046 5694 436102
rect 5762 436046 5818 436102
rect 5886 436046 5942 436102
rect 5514 435922 5570 435978
rect 5638 435922 5694 435978
rect 5762 435922 5818 435978
rect 5886 435922 5942 435978
rect -860 418294 -804 418350
rect -736 418294 -680 418350
rect -612 418294 -556 418350
rect -488 418294 -432 418350
rect -860 418170 -804 418226
rect -736 418170 -680 418226
rect -612 418170 -556 418226
rect -488 418170 -432 418226
rect -860 418046 -804 418102
rect -736 418046 -680 418102
rect -612 418046 -556 418102
rect -488 418046 -432 418102
rect -860 417922 -804 417978
rect -736 417922 -680 417978
rect -612 417922 -556 417978
rect -488 417922 -432 417978
rect 12518 436294 12574 436350
rect 12642 436294 12698 436350
rect 12518 436170 12574 436226
rect 12642 436170 12698 436226
rect 12518 436046 12574 436102
rect 12642 436046 12698 436102
rect 12518 435922 12574 435978
rect 12642 435922 12698 435978
rect 43238 436294 43294 436350
rect 43362 436294 43418 436350
rect 43238 436170 43294 436226
rect 43362 436170 43418 436226
rect 43238 436046 43294 436102
rect 43362 436046 43418 436102
rect 43238 435922 43294 435978
rect 43362 435922 43418 435978
rect 73958 436294 74014 436350
rect 74082 436294 74138 436350
rect 73958 436170 74014 436226
rect 74082 436170 74138 436226
rect 73958 436046 74014 436102
rect 74082 436046 74138 436102
rect 73958 435922 74014 435978
rect 74082 435922 74138 435978
rect 104678 436294 104734 436350
rect 104802 436294 104858 436350
rect 104678 436170 104734 436226
rect 104802 436170 104858 436226
rect 104678 436046 104734 436102
rect 104802 436046 104858 436102
rect 104678 435922 104734 435978
rect 104802 435922 104858 435978
rect 135398 436294 135454 436350
rect 135522 436294 135578 436350
rect 135398 436170 135454 436226
rect 135522 436170 135578 436226
rect 135398 436046 135454 436102
rect 135522 436046 135578 436102
rect 135398 435922 135454 435978
rect 135522 435922 135578 435978
rect 166118 436294 166174 436350
rect 166242 436294 166298 436350
rect 166118 436170 166174 436226
rect 166242 436170 166298 436226
rect 166118 436046 166174 436102
rect 166242 436046 166298 436102
rect 166118 435922 166174 435978
rect 166242 435922 166298 435978
rect 196838 436294 196894 436350
rect 196962 436294 197018 436350
rect 196838 436170 196894 436226
rect 196962 436170 197018 436226
rect 196838 436046 196894 436102
rect 196962 436046 197018 436102
rect 196838 435922 196894 435978
rect 196962 435922 197018 435978
rect 227558 436294 227614 436350
rect 227682 436294 227738 436350
rect 227558 436170 227614 436226
rect 227682 436170 227738 436226
rect 227558 436046 227614 436102
rect 227682 436046 227738 436102
rect 227558 435922 227614 435978
rect 227682 435922 227738 435978
rect 258278 436294 258334 436350
rect 258402 436294 258458 436350
rect 258278 436170 258334 436226
rect 258402 436170 258458 436226
rect 258278 436046 258334 436102
rect 258402 436046 258458 436102
rect 258278 435922 258334 435978
rect 258402 435922 258458 435978
rect 288998 436294 289054 436350
rect 289122 436294 289178 436350
rect 288998 436170 289054 436226
rect 289122 436170 289178 436226
rect 288998 436046 289054 436102
rect 289122 436046 289178 436102
rect 288998 435922 289054 435978
rect 289122 435922 289178 435978
rect 319718 436294 319774 436350
rect 319842 436294 319898 436350
rect 319718 436170 319774 436226
rect 319842 436170 319898 436226
rect 319718 436046 319774 436102
rect 319842 436046 319898 436102
rect 319718 435922 319774 435978
rect 319842 435922 319898 435978
rect 350438 436294 350494 436350
rect 350562 436294 350618 436350
rect 350438 436170 350494 436226
rect 350562 436170 350618 436226
rect 350438 436046 350494 436102
rect 350562 436046 350618 436102
rect 350438 435922 350494 435978
rect 350562 435922 350618 435978
rect 381158 436294 381214 436350
rect 381282 436294 381338 436350
rect 381158 436170 381214 436226
rect 381282 436170 381338 436226
rect 381158 436046 381214 436102
rect 381282 436046 381338 436102
rect 381158 435922 381214 435978
rect 381282 435922 381338 435978
rect 411878 436294 411934 436350
rect 412002 436294 412058 436350
rect 411878 436170 411934 436226
rect 412002 436170 412058 436226
rect 411878 436046 411934 436102
rect 412002 436046 412058 436102
rect 411878 435922 411934 435978
rect 412002 435922 412058 435978
rect 442598 436294 442654 436350
rect 442722 436294 442778 436350
rect 442598 436170 442654 436226
rect 442722 436170 442778 436226
rect 442598 436046 442654 436102
rect 442722 436046 442778 436102
rect 442598 435922 442654 435978
rect 442722 435922 442778 435978
rect 473318 436294 473374 436350
rect 473442 436294 473498 436350
rect 473318 436170 473374 436226
rect 473442 436170 473498 436226
rect 473318 436046 473374 436102
rect 473442 436046 473498 436102
rect 473318 435922 473374 435978
rect 473442 435922 473498 435978
rect 504038 436294 504094 436350
rect 504162 436294 504218 436350
rect 504038 436170 504094 436226
rect 504162 436170 504218 436226
rect 504038 436046 504094 436102
rect 504162 436046 504218 436102
rect 504038 435922 504094 435978
rect 504162 435922 504218 435978
rect 534758 436294 534814 436350
rect 534882 436294 534938 436350
rect 534758 436170 534814 436226
rect 534882 436170 534938 436226
rect 534758 436046 534814 436102
rect 534882 436046 534938 436102
rect 534758 435922 534814 435978
rect 534882 435922 534938 435978
rect 565478 436294 565534 436350
rect 565602 436294 565658 436350
rect 565478 436170 565534 436226
rect 565602 436170 565658 436226
rect 565478 436046 565534 436102
rect 565602 436046 565658 436102
rect 565478 435922 565534 435978
rect 565602 435922 565658 435978
rect 592914 460294 592970 460350
rect 593038 460294 593094 460350
rect 593162 460294 593218 460350
rect 593286 460294 593342 460350
rect 592914 460170 592970 460226
rect 593038 460170 593094 460226
rect 593162 460170 593218 460226
rect 593286 460170 593342 460226
rect 592914 460046 592970 460102
rect 593038 460046 593094 460102
rect 593162 460046 593218 460102
rect 593286 460046 593342 460102
rect 592914 459922 592970 459978
rect 593038 459922 593094 459978
rect 593162 459922 593218 459978
rect 593286 459922 593342 459978
rect 589194 436294 589250 436350
rect 589318 436294 589374 436350
rect 589442 436294 589498 436350
rect 589566 436294 589622 436350
rect 589194 436170 589250 436226
rect 589318 436170 589374 436226
rect 589442 436170 589498 436226
rect 589566 436170 589622 436226
rect 589194 436046 589250 436102
rect 589318 436046 589374 436102
rect 589442 436046 589498 436102
rect 589566 436046 589622 436102
rect 589194 435922 589250 435978
rect 589318 435922 589374 435978
rect 589442 435922 589498 435978
rect 589566 435922 589622 435978
rect 5514 418294 5570 418350
rect 5638 418294 5694 418350
rect 5762 418294 5818 418350
rect 5886 418294 5942 418350
rect 5514 418170 5570 418226
rect 5638 418170 5694 418226
rect 5762 418170 5818 418226
rect 5886 418170 5942 418226
rect 5514 418046 5570 418102
rect 5638 418046 5694 418102
rect 5762 418046 5818 418102
rect 5886 418046 5942 418102
rect 5514 417922 5570 417978
rect 5638 417922 5694 417978
rect 5762 417922 5818 417978
rect 5886 417922 5942 417978
rect -860 400294 -804 400350
rect -736 400294 -680 400350
rect -612 400294 -556 400350
rect -488 400294 -432 400350
rect -860 400170 -804 400226
rect -736 400170 -680 400226
rect -612 400170 -556 400226
rect -488 400170 -432 400226
rect -860 400046 -804 400102
rect -736 400046 -680 400102
rect -612 400046 -556 400102
rect -488 400046 -432 400102
rect -860 399922 -804 399978
rect -736 399922 -680 399978
rect -612 399922 -556 399978
rect -488 399922 -432 399978
rect 5514 400294 5570 400350
rect 5638 400294 5694 400350
rect 5762 400294 5818 400350
rect 5886 400294 5942 400350
rect 5514 400170 5570 400226
rect 5638 400170 5694 400226
rect 5762 400170 5818 400226
rect 5886 400170 5942 400226
rect 5514 400046 5570 400102
rect 5638 400046 5694 400102
rect 5762 400046 5818 400102
rect 5886 400046 5942 400102
rect 5514 399922 5570 399978
rect 5638 399922 5694 399978
rect 5762 399922 5818 399978
rect 5886 399922 5942 399978
rect -860 382294 -804 382350
rect -736 382294 -680 382350
rect -612 382294 -556 382350
rect -488 382294 -432 382350
rect -860 382170 -804 382226
rect -736 382170 -680 382226
rect -612 382170 -556 382226
rect -488 382170 -432 382226
rect -860 382046 -804 382102
rect -736 382046 -680 382102
rect -612 382046 -556 382102
rect -488 382046 -432 382102
rect -860 381922 -804 381978
rect -736 381922 -680 381978
rect -612 381922 -556 381978
rect -488 381922 -432 381978
rect -860 364294 -804 364350
rect -736 364294 -680 364350
rect -612 364294 -556 364350
rect -488 364294 -432 364350
rect -860 364170 -804 364226
rect -736 364170 -680 364226
rect -612 364170 -556 364226
rect -488 364170 -432 364226
rect -860 364046 -804 364102
rect -736 364046 -680 364102
rect -612 364046 -556 364102
rect -488 364046 -432 364102
rect -860 363922 -804 363978
rect -736 363922 -680 363978
rect -612 363922 -556 363978
rect -488 363922 -432 363978
rect 27878 424294 27934 424350
rect 28002 424294 28058 424350
rect 27878 424170 27934 424226
rect 28002 424170 28058 424226
rect 27878 424046 27934 424102
rect 28002 424046 28058 424102
rect 27878 423922 27934 423978
rect 28002 423922 28058 423978
rect 58598 424294 58654 424350
rect 58722 424294 58778 424350
rect 58598 424170 58654 424226
rect 58722 424170 58778 424226
rect 58598 424046 58654 424102
rect 58722 424046 58778 424102
rect 58598 423922 58654 423978
rect 58722 423922 58778 423978
rect 89318 424294 89374 424350
rect 89442 424294 89498 424350
rect 89318 424170 89374 424226
rect 89442 424170 89498 424226
rect 89318 424046 89374 424102
rect 89442 424046 89498 424102
rect 89318 423922 89374 423978
rect 89442 423922 89498 423978
rect 120038 424294 120094 424350
rect 120162 424294 120218 424350
rect 120038 424170 120094 424226
rect 120162 424170 120218 424226
rect 120038 424046 120094 424102
rect 120162 424046 120218 424102
rect 120038 423922 120094 423978
rect 120162 423922 120218 423978
rect 150758 424294 150814 424350
rect 150882 424294 150938 424350
rect 150758 424170 150814 424226
rect 150882 424170 150938 424226
rect 150758 424046 150814 424102
rect 150882 424046 150938 424102
rect 150758 423922 150814 423978
rect 150882 423922 150938 423978
rect 181478 424294 181534 424350
rect 181602 424294 181658 424350
rect 181478 424170 181534 424226
rect 181602 424170 181658 424226
rect 181478 424046 181534 424102
rect 181602 424046 181658 424102
rect 181478 423922 181534 423978
rect 181602 423922 181658 423978
rect 212198 424294 212254 424350
rect 212322 424294 212378 424350
rect 212198 424170 212254 424226
rect 212322 424170 212378 424226
rect 212198 424046 212254 424102
rect 212322 424046 212378 424102
rect 212198 423922 212254 423978
rect 212322 423922 212378 423978
rect 242918 424294 242974 424350
rect 243042 424294 243098 424350
rect 242918 424170 242974 424226
rect 243042 424170 243098 424226
rect 242918 424046 242974 424102
rect 243042 424046 243098 424102
rect 242918 423922 242974 423978
rect 243042 423922 243098 423978
rect 273638 424294 273694 424350
rect 273762 424294 273818 424350
rect 273638 424170 273694 424226
rect 273762 424170 273818 424226
rect 273638 424046 273694 424102
rect 273762 424046 273818 424102
rect 273638 423922 273694 423978
rect 273762 423922 273818 423978
rect 304358 424294 304414 424350
rect 304482 424294 304538 424350
rect 304358 424170 304414 424226
rect 304482 424170 304538 424226
rect 304358 424046 304414 424102
rect 304482 424046 304538 424102
rect 304358 423922 304414 423978
rect 304482 423922 304538 423978
rect 335078 424294 335134 424350
rect 335202 424294 335258 424350
rect 335078 424170 335134 424226
rect 335202 424170 335258 424226
rect 335078 424046 335134 424102
rect 335202 424046 335258 424102
rect 335078 423922 335134 423978
rect 335202 423922 335258 423978
rect 365798 424294 365854 424350
rect 365922 424294 365978 424350
rect 365798 424170 365854 424226
rect 365922 424170 365978 424226
rect 365798 424046 365854 424102
rect 365922 424046 365978 424102
rect 365798 423922 365854 423978
rect 365922 423922 365978 423978
rect 396518 424294 396574 424350
rect 396642 424294 396698 424350
rect 396518 424170 396574 424226
rect 396642 424170 396698 424226
rect 396518 424046 396574 424102
rect 396642 424046 396698 424102
rect 396518 423922 396574 423978
rect 396642 423922 396698 423978
rect 427238 424294 427294 424350
rect 427362 424294 427418 424350
rect 427238 424170 427294 424226
rect 427362 424170 427418 424226
rect 427238 424046 427294 424102
rect 427362 424046 427418 424102
rect 427238 423922 427294 423978
rect 427362 423922 427418 423978
rect 457958 424294 458014 424350
rect 458082 424294 458138 424350
rect 457958 424170 458014 424226
rect 458082 424170 458138 424226
rect 457958 424046 458014 424102
rect 458082 424046 458138 424102
rect 457958 423922 458014 423978
rect 458082 423922 458138 423978
rect 488678 424294 488734 424350
rect 488802 424294 488858 424350
rect 488678 424170 488734 424226
rect 488802 424170 488858 424226
rect 488678 424046 488734 424102
rect 488802 424046 488858 424102
rect 488678 423922 488734 423978
rect 488802 423922 488858 423978
rect 519398 424294 519454 424350
rect 519522 424294 519578 424350
rect 519398 424170 519454 424226
rect 519522 424170 519578 424226
rect 519398 424046 519454 424102
rect 519522 424046 519578 424102
rect 519398 423922 519454 423978
rect 519522 423922 519578 423978
rect 550118 424294 550174 424350
rect 550242 424294 550298 424350
rect 550118 424170 550174 424226
rect 550242 424170 550298 424226
rect 550118 424046 550174 424102
rect 550242 424046 550298 424102
rect 550118 423922 550174 423978
rect 550242 423922 550298 423978
rect 12518 418294 12574 418350
rect 12642 418294 12698 418350
rect 12518 418170 12574 418226
rect 12642 418170 12698 418226
rect 12518 418046 12574 418102
rect 12642 418046 12698 418102
rect 12518 417922 12574 417978
rect 12642 417922 12698 417978
rect 43238 418294 43294 418350
rect 43362 418294 43418 418350
rect 43238 418170 43294 418226
rect 43362 418170 43418 418226
rect 43238 418046 43294 418102
rect 43362 418046 43418 418102
rect 43238 417922 43294 417978
rect 43362 417922 43418 417978
rect 73958 418294 74014 418350
rect 74082 418294 74138 418350
rect 73958 418170 74014 418226
rect 74082 418170 74138 418226
rect 73958 418046 74014 418102
rect 74082 418046 74138 418102
rect 73958 417922 74014 417978
rect 74082 417922 74138 417978
rect 104678 418294 104734 418350
rect 104802 418294 104858 418350
rect 104678 418170 104734 418226
rect 104802 418170 104858 418226
rect 104678 418046 104734 418102
rect 104802 418046 104858 418102
rect 104678 417922 104734 417978
rect 104802 417922 104858 417978
rect 135398 418294 135454 418350
rect 135522 418294 135578 418350
rect 135398 418170 135454 418226
rect 135522 418170 135578 418226
rect 135398 418046 135454 418102
rect 135522 418046 135578 418102
rect 135398 417922 135454 417978
rect 135522 417922 135578 417978
rect 166118 418294 166174 418350
rect 166242 418294 166298 418350
rect 166118 418170 166174 418226
rect 166242 418170 166298 418226
rect 166118 418046 166174 418102
rect 166242 418046 166298 418102
rect 166118 417922 166174 417978
rect 166242 417922 166298 417978
rect 196838 418294 196894 418350
rect 196962 418294 197018 418350
rect 196838 418170 196894 418226
rect 196962 418170 197018 418226
rect 196838 418046 196894 418102
rect 196962 418046 197018 418102
rect 196838 417922 196894 417978
rect 196962 417922 197018 417978
rect 227558 418294 227614 418350
rect 227682 418294 227738 418350
rect 227558 418170 227614 418226
rect 227682 418170 227738 418226
rect 227558 418046 227614 418102
rect 227682 418046 227738 418102
rect 227558 417922 227614 417978
rect 227682 417922 227738 417978
rect 258278 418294 258334 418350
rect 258402 418294 258458 418350
rect 258278 418170 258334 418226
rect 258402 418170 258458 418226
rect 258278 418046 258334 418102
rect 258402 418046 258458 418102
rect 258278 417922 258334 417978
rect 258402 417922 258458 417978
rect 288998 418294 289054 418350
rect 289122 418294 289178 418350
rect 288998 418170 289054 418226
rect 289122 418170 289178 418226
rect 288998 418046 289054 418102
rect 289122 418046 289178 418102
rect 288998 417922 289054 417978
rect 289122 417922 289178 417978
rect 319718 418294 319774 418350
rect 319842 418294 319898 418350
rect 319718 418170 319774 418226
rect 319842 418170 319898 418226
rect 319718 418046 319774 418102
rect 319842 418046 319898 418102
rect 319718 417922 319774 417978
rect 319842 417922 319898 417978
rect 350438 418294 350494 418350
rect 350562 418294 350618 418350
rect 350438 418170 350494 418226
rect 350562 418170 350618 418226
rect 350438 418046 350494 418102
rect 350562 418046 350618 418102
rect 350438 417922 350494 417978
rect 350562 417922 350618 417978
rect 381158 418294 381214 418350
rect 381282 418294 381338 418350
rect 381158 418170 381214 418226
rect 381282 418170 381338 418226
rect 381158 418046 381214 418102
rect 381282 418046 381338 418102
rect 381158 417922 381214 417978
rect 381282 417922 381338 417978
rect 411878 418294 411934 418350
rect 412002 418294 412058 418350
rect 411878 418170 411934 418226
rect 412002 418170 412058 418226
rect 411878 418046 411934 418102
rect 412002 418046 412058 418102
rect 411878 417922 411934 417978
rect 412002 417922 412058 417978
rect 442598 418294 442654 418350
rect 442722 418294 442778 418350
rect 442598 418170 442654 418226
rect 442722 418170 442778 418226
rect 442598 418046 442654 418102
rect 442722 418046 442778 418102
rect 442598 417922 442654 417978
rect 442722 417922 442778 417978
rect 473318 418294 473374 418350
rect 473442 418294 473498 418350
rect 473318 418170 473374 418226
rect 473442 418170 473498 418226
rect 473318 418046 473374 418102
rect 473442 418046 473498 418102
rect 473318 417922 473374 417978
rect 473442 417922 473498 417978
rect 504038 418294 504094 418350
rect 504162 418294 504218 418350
rect 504038 418170 504094 418226
rect 504162 418170 504218 418226
rect 504038 418046 504094 418102
rect 504162 418046 504218 418102
rect 504038 417922 504094 417978
rect 504162 417922 504218 417978
rect 534758 418294 534814 418350
rect 534882 418294 534938 418350
rect 534758 418170 534814 418226
rect 534882 418170 534938 418226
rect 534758 418046 534814 418102
rect 534882 418046 534938 418102
rect 534758 417922 534814 417978
rect 534882 417922 534938 417978
rect 565478 418294 565534 418350
rect 565602 418294 565658 418350
rect 565478 418170 565534 418226
rect 565602 418170 565658 418226
rect 565478 418046 565534 418102
rect 565602 418046 565658 418102
rect 565478 417922 565534 417978
rect 565602 417922 565658 417978
rect 27878 406294 27934 406350
rect 28002 406294 28058 406350
rect 27878 406170 27934 406226
rect 28002 406170 28058 406226
rect 27878 406046 27934 406102
rect 28002 406046 28058 406102
rect 27878 405922 27934 405978
rect 28002 405922 28058 405978
rect 58598 406294 58654 406350
rect 58722 406294 58778 406350
rect 58598 406170 58654 406226
rect 58722 406170 58778 406226
rect 58598 406046 58654 406102
rect 58722 406046 58778 406102
rect 58598 405922 58654 405978
rect 58722 405922 58778 405978
rect 89318 406294 89374 406350
rect 89442 406294 89498 406350
rect 89318 406170 89374 406226
rect 89442 406170 89498 406226
rect 89318 406046 89374 406102
rect 89442 406046 89498 406102
rect 89318 405922 89374 405978
rect 89442 405922 89498 405978
rect 120038 406294 120094 406350
rect 120162 406294 120218 406350
rect 120038 406170 120094 406226
rect 120162 406170 120218 406226
rect 120038 406046 120094 406102
rect 120162 406046 120218 406102
rect 120038 405922 120094 405978
rect 120162 405922 120218 405978
rect 150758 406294 150814 406350
rect 150882 406294 150938 406350
rect 150758 406170 150814 406226
rect 150882 406170 150938 406226
rect 150758 406046 150814 406102
rect 150882 406046 150938 406102
rect 150758 405922 150814 405978
rect 150882 405922 150938 405978
rect 181478 406294 181534 406350
rect 181602 406294 181658 406350
rect 181478 406170 181534 406226
rect 181602 406170 181658 406226
rect 181478 406046 181534 406102
rect 181602 406046 181658 406102
rect 181478 405922 181534 405978
rect 181602 405922 181658 405978
rect 212198 406294 212254 406350
rect 212322 406294 212378 406350
rect 212198 406170 212254 406226
rect 212322 406170 212378 406226
rect 212198 406046 212254 406102
rect 212322 406046 212378 406102
rect 212198 405922 212254 405978
rect 212322 405922 212378 405978
rect 242918 406294 242974 406350
rect 243042 406294 243098 406350
rect 242918 406170 242974 406226
rect 243042 406170 243098 406226
rect 242918 406046 242974 406102
rect 243042 406046 243098 406102
rect 242918 405922 242974 405978
rect 243042 405922 243098 405978
rect 273638 406294 273694 406350
rect 273762 406294 273818 406350
rect 273638 406170 273694 406226
rect 273762 406170 273818 406226
rect 273638 406046 273694 406102
rect 273762 406046 273818 406102
rect 273638 405922 273694 405978
rect 273762 405922 273818 405978
rect 304358 406294 304414 406350
rect 304482 406294 304538 406350
rect 304358 406170 304414 406226
rect 304482 406170 304538 406226
rect 304358 406046 304414 406102
rect 304482 406046 304538 406102
rect 304358 405922 304414 405978
rect 304482 405922 304538 405978
rect 335078 406294 335134 406350
rect 335202 406294 335258 406350
rect 335078 406170 335134 406226
rect 335202 406170 335258 406226
rect 335078 406046 335134 406102
rect 335202 406046 335258 406102
rect 335078 405922 335134 405978
rect 335202 405922 335258 405978
rect 365798 406294 365854 406350
rect 365922 406294 365978 406350
rect 365798 406170 365854 406226
rect 365922 406170 365978 406226
rect 365798 406046 365854 406102
rect 365922 406046 365978 406102
rect 365798 405922 365854 405978
rect 365922 405922 365978 405978
rect 396518 406294 396574 406350
rect 396642 406294 396698 406350
rect 396518 406170 396574 406226
rect 396642 406170 396698 406226
rect 396518 406046 396574 406102
rect 396642 406046 396698 406102
rect 396518 405922 396574 405978
rect 396642 405922 396698 405978
rect 427238 406294 427294 406350
rect 427362 406294 427418 406350
rect 427238 406170 427294 406226
rect 427362 406170 427418 406226
rect 427238 406046 427294 406102
rect 427362 406046 427418 406102
rect 427238 405922 427294 405978
rect 427362 405922 427418 405978
rect 457958 406294 458014 406350
rect 458082 406294 458138 406350
rect 457958 406170 458014 406226
rect 458082 406170 458138 406226
rect 457958 406046 458014 406102
rect 458082 406046 458138 406102
rect 457958 405922 458014 405978
rect 458082 405922 458138 405978
rect 488678 406294 488734 406350
rect 488802 406294 488858 406350
rect 488678 406170 488734 406226
rect 488802 406170 488858 406226
rect 488678 406046 488734 406102
rect 488802 406046 488858 406102
rect 488678 405922 488734 405978
rect 488802 405922 488858 405978
rect 519398 406294 519454 406350
rect 519522 406294 519578 406350
rect 519398 406170 519454 406226
rect 519522 406170 519578 406226
rect 519398 406046 519454 406102
rect 519522 406046 519578 406102
rect 519398 405922 519454 405978
rect 519522 405922 519578 405978
rect 550118 406294 550174 406350
rect 550242 406294 550298 406350
rect 550118 406170 550174 406226
rect 550242 406170 550298 406226
rect 550118 406046 550174 406102
rect 550242 406046 550298 406102
rect 550118 405922 550174 405978
rect 550242 405922 550298 405978
rect 592914 442294 592970 442350
rect 593038 442294 593094 442350
rect 593162 442294 593218 442350
rect 593286 442294 593342 442350
rect 592914 442170 592970 442226
rect 593038 442170 593094 442226
rect 593162 442170 593218 442226
rect 593286 442170 593342 442226
rect 592914 442046 592970 442102
rect 593038 442046 593094 442102
rect 593162 442046 593218 442102
rect 593286 442046 593342 442102
rect 592914 441922 592970 441978
rect 593038 441922 593094 441978
rect 593162 441922 593218 441978
rect 593286 441922 593342 441978
rect 589194 418294 589250 418350
rect 589318 418294 589374 418350
rect 589442 418294 589498 418350
rect 589566 418294 589622 418350
rect 589194 418170 589250 418226
rect 589318 418170 589374 418226
rect 589442 418170 589498 418226
rect 589566 418170 589622 418226
rect 589194 418046 589250 418102
rect 589318 418046 589374 418102
rect 589442 418046 589498 418102
rect 589566 418046 589622 418102
rect 589194 417922 589250 417978
rect 589318 417922 589374 417978
rect 589442 417922 589498 417978
rect 589566 417922 589622 417978
rect 12518 400294 12574 400350
rect 12642 400294 12698 400350
rect 12518 400170 12574 400226
rect 12642 400170 12698 400226
rect 12518 400046 12574 400102
rect 12642 400046 12698 400102
rect 12518 399922 12574 399978
rect 12642 399922 12698 399978
rect 43238 400294 43294 400350
rect 43362 400294 43418 400350
rect 43238 400170 43294 400226
rect 43362 400170 43418 400226
rect 43238 400046 43294 400102
rect 43362 400046 43418 400102
rect 43238 399922 43294 399978
rect 43362 399922 43418 399978
rect 73958 400294 74014 400350
rect 74082 400294 74138 400350
rect 73958 400170 74014 400226
rect 74082 400170 74138 400226
rect 73958 400046 74014 400102
rect 74082 400046 74138 400102
rect 73958 399922 74014 399978
rect 74082 399922 74138 399978
rect 104678 400294 104734 400350
rect 104802 400294 104858 400350
rect 104678 400170 104734 400226
rect 104802 400170 104858 400226
rect 104678 400046 104734 400102
rect 104802 400046 104858 400102
rect 104678 399922 104734 399978
rect 104802 399922 104858 399978
rect 135398 400294 135454 400350
rect 135522 400294 135578 400350
rect 135398 400170 135454 400226
rect 135522 400170 135578 400226
rect 135398 400046 135454 400102
rect 135522 400046 135578 400102
rect 135398 399922 135454 399978
rect 135522 399922 135578 399978
rect 166118 400294 166174 400350
rect 166242 400294 166298 400350
rect 166118 400170 166174 400226
rect 166242 400170 166298 400226
rect 166118 400046 166174 400102
rect 166242 400046 166298 400102
rect 166118 399922 166174 399978
rect 166242 399922 166298 399978
rect 196838 400294 196894 400350
rect 196962 400294 197018 400350
rect 196838 400170 196894 400226
rect 196962 400170 197018 400226
rect 196838 400046 196894 400102
rect 196962 400046 197018 400102
rect 196838 399922 196894 399978
rect 196962 399922 197018 399978
rect 227558 400294 227614 400350
rect 227682 400294 227738 400350
rect 227558 400170 227614 400226
rect 227682 400170 227738 400226
rect 227558 400046 227614 400102
rect 227682 400046 227738 400102
rect 227558 399922 227614 399978
rect 227682 399922 227738 399978
rect 258278 400294 258334 400350
rect 258402 400294 258458 400350
rect 258278 400170 258334 400226
rect 258402 400170 258458 400226
rect 258278 400046 258334 400102
rect 258402 400046 258458 400102
rect 258278 399922 258334 399978
rect 258402 399922 258458 399978
rect 288998 400294 289054 400350
rect 289122 400294 289178 400350
rect 288998 400170 289054 400226
rect 289122 400170 289178 400226
rect 288998 400046 289054 400102
rect 289122 400046 289178 400102
rect 288998 399922 289054 399978
rect 289122 399922 289178 399978
rect 319718 400294 319774 400350
rect 319842 400294 319898 400350
rect 319718 400170 319774 400226
rect 319842 400170 319898 400226
rect 319718 400046 319774 400102
rect 319842 400046 319898 400102
rect 319718 399922 319774 399978
rect 319842 399922 319898 399978
rect 350438 400294 350494 400350
rect 350562 400294 350618 400350
rect 350438 400170 350494 400226
rect 350562 400170 350618 400226
rect 350438 400046 350494 400102
rect 350562 400046 350618 400102
rect 350438 399922 350494 399978
rect 350562 399922 350618 399978
rect 381158 400294 381214 400350
rect 381282 400294 381338 400350
rect 381158 400170 381214 400226
rect 381282 400170 381338 400226
rect 381158 400046 381214 400102
rect 381282 400046 381338 400102
rect 381158 399922 381214 399978
rect 381282 399922 381338 399978
rect 411878 400294 411934 400350
rect 412002 400294 412058 400350
rect 411878 400170 411934 400226
rect 412002 400170 412058 400226
rect 411878 400046 411934 400102
rect 412002 400046 412058 400102
rect 411878 399922 411934 399978
rect 412002 399922 412058 399978
rect 442598 400294 442654 400350
rect 442722 400294 442778 400350
rect 442598 400170 442654 400226
rect 442722 400170 442778 400226
rect 442598 400046 442654 400102
rect 442722 400046 442778 400102
rect 442598 399922 442654 399978
rect 442722 399922 442778 399978
rect 473318 400294 473374 400350
rect 473442 400294 473498 400350
rect 473318 400170 473374 400226
rect 473442 400170 473498 400226
rect 473318 400046 473374 400102
rect 473442 400046 473498 400102
rect 473318 399922 473374 399978
rect 473442 399922 473498 399978
rect 504038 400294 504094 400350
rect 504162 400294 504218 400350
rect 504038 400170 504094 400226
rect 504162 400170 504218 400226
rect 504038 400046 504094 400102
rect 504162 400046 504218 400102
rect 504038 399922 504094 399978
rect 504162 399922 504218 399978
rect 534758 400294 534814 400350
rect 534882 400294 534938 400350
rect 534758 400170 534814 400226
rect 534882 400170 534938 400226
rect 534758 400046 534814 400102
rect 534882 400046 534938 400102
rect 534758 399922 534814 399978
rect 534882 399922 534938 399978
rect 565478 400294 565534 400350
rect 565602 400294 565658 400350
rect 565478 400170 565534 400226
rect 565602 400170 565658 400226
rect 565478 400046 565534 400102
rect 565602 400046 565658 400102
rect 565478 399922 565534 399978
rect 565602 399922 565658 399978
rect 5514 382294 5570 382350
rect 5638 382294 5694 382350
rect 5762 382294 5818 382350
rect 5886 382294 5942 382350
rect 5514 382170 5570 382226
rect 5638 382170 5694 382226
rect 5762 382170 5818 382226
rect 5886 382170 5942 382226
rect 5514 382046 5570 382102
rect 5638 382046 5694 382102
rect 5762 382046 5818 382102
rect 5886 382046 5942 382102
rect 5514 381922 5570 381978
rect 5638 381922 5694 381978
rect 5762 381922 5818 381978
rect 5886 381922 5942 381978
rect 27878 388294 27934 388350
rect 28002 388294 28058 388350
rect 27878 388170 27934 388226
rect 28002 388170 28058 388226
rect 27878 388046 27934 388102
rect 28002 388046 28058 388102
rect 27878 387922 27934 387978
rect 28002 387922 28058 387978
rect 58598 388294 58654 388350
rect 58722 388294 58778 388350
rect 58598 388170 58654 388226
rect 58722 388170 58778 388226
rect 58598 388046 58654 388102
rect 58722 388046 58778 388102
rect 58598 387922 58654 387978
rect 58722 387922 58778 387978
rect 89318 388294 89374 388350
rect 89442 388294 89498 388350
rect 89318 388170 89374 388226
rect 89442 388170 89498 388226
rect 89318 388046 89374 388102
rect 89442 388046 89498 388102
rect 89318 387922 89374 387978
rect 89442 387922 89498 387978
rect 120038 388294 120094 388350
rect 120162 388294 120218 388350
rect 120038 388170 120094 388226
rect 120162 388170 120218 388226
rect 120038 388046 120094 388102
rect 120162 388046 120218 388102
rect 120038 387922 120094 387978
rect 120162 387922 120218 387978
rect 150758 388294 150814 388350
rect 150882 388294 150938 388350
rect 150758 388170 150814 388226
rect 150882 388170 150938 388226
rect 150758 388046 150814 388102
rect 150882 388046 150938 388102
rect 150758 387922 150814 387978
rect 150882 387922 150938 387978
rect 181478 388294 181534 388350
rect 181602 388294 181658 388350
rect 181478 388170 181534 388226
rect 181602 388170 181658 388226
rect 181478 388046 181534 388102
rect 181602 388046 181658 388102
rect 181478 387922 181534 387978
rect 181602 387922 181658 387978
rect 212198 388294 212254 388350
rect 212322 388294 212378 388350
rect 212198 388170 212254 388226
rect 212322 388170 212378 388226
rect 212198 388046 212254 388102
rect 212322 388046 212378 388102
rect 212198 387922 212254 387978
rect 212322 387922 212378 387978
rect 242918 388294 242974 388350
rect 243042 388294 243098 388350
rect 242918 388170 242974 388226
rect 243042 388170 243098 388226
rect 242918 388046 242974 388102
rect 243042 388046 243098 388102
rect 242918 387922 242974 387978
rect 243042 387922 243098 387978
rect 273638 388294 273694 388350
rect 273762 388294 273818 388350
rect 273638 388170 273694 388226
rect 273762 388170 273818 388226
rect 273638 388046 273694 388102
rect 273762 388046 273818 388102
rect 273638 387922 273694 387978
rect 273762 387922 273818 387978
rect 304358 388294 304414 388350
rect 304482 388294 304538 388350
rect 304358 388170 304414 388226
rect 304482 388170 304538 388226
rect 304358 388046 304414 388102
rect 304482 388046 304538 388102
rect 304358 387922 304414 387978
rect 304482 387922 304538 387978
rect 335078 388294 335134 388350
rect 335202 388294 335258 388350
rect 335078 388170 335134 388226
rect 335202 388170 335258 388226
rect 335078 388046 335134 388102
rect 335202 388046 335258 388102
rect 335078 387922 335134 387978
rect 335202 387922 335258 387978
rect 365798 388294 365854 388350
rect 365922 388294 365978 388350
rect 365798 388170 365854 388226
rect 365922 388170 365978 388226
rect 365798 388046 365854 388102
rect 365922 388046 365978 388102
rect 365798 387922 365854 387978
rect 365922 387922 365978 387978
rect 396518 388294 396574 388350
rect 396642 388294 396698 388350
rect 396518 388170 396574 388226
rect 396642 388170 396698 388226
rect 396518 388046 396574 388102
rect 396642 388046 396698 388102
rect 396518 387922 396574 387978
rect 396642 387922 396698 387978
rect 427238 388294 427294 388350
rect 427362 388294 427418 388350
rect 427238 388170 427294 388226
rect 427362 388170 427418 388226
rect 427238 388046 427294 388102
rect 427362 388046 427418 388102
rect 427238 387922 427294 387978
rect 427362 387922 427418 387978
rect 457958 388294 458014 388350
rect 458082 388294 458138 388350
rect 457958 388170 458014 388226
rect 458082 388170 458138 388226
rect 457958 388046 458014 388102
rect 458082 388046 458138 388102
rect 457958 387922 458014 387978
rect 458082 387922 458138 387978
rect 488678 388294 488734 388350
rect 488802 388294 488858 388350
rect 488678 388170 488734 388226
rect 488802 388170 488858 388226
rect 488678 388046 488734 388102
rect 488802 388046 488858 388102
rect 488678 387922 488734 387978
rect 488802 387922 488858 387978
rect 519398 388294 519454 388350
rect 519522 388294 519578 388350
rect 519398 388170 519454 388226
rect 519522 388170 519578 388226
rect 519398 388046 519454 388102
rect 519522 388046 519578 388102
rect 519398 387922 519454 387978
rect 519522 387922 519578 387978
rect 550118 388294 550174 388350
rect 550242 388294 550298 388350
rect 550118 388170 550174 388226
rect 550242 388170 550298 388226
rect 550118 388046 550174 388102
rect 550242 388046 550298 388102
rect 550118 387922 550174 387978
rect 550242 387922 550298 387978
rect 12518 382294 12574 382350
rect 12642 382294 12698 382350
rect 12518 382170 12574 382226
rect 12642 382170 12698 382226
rect 12518 382046 12574 382102
rect 12642 382046 12698 382102
rect 12518 381922 12574 381978
rect 12642 381922 12698 381978
rect 43238 382294 43294 382350
rect 43362 382294 43418 382350
rect 43238 382170 43294 382226
rect 43362 382170 43418 382226
rect 43238 382046 43294 382102
rect 43362 382046 43418 382102
rect 43238 381922 43294 381978
rect 43362 381922 43418 381978
rect 73958 382294 74014 382350
rect 74082 382294 74138 382350
rect 73958 382170 74014 382226
rect 74082 382170 74138 382226
rect 73958 382046 74014 382102
rect 74082 382046 74138 382102
rect 73958 381922 74014 381978
rect 74082 381922 74138 381978
rect 104678 382294 104734 382350
rect 104802 382294 104858 382350
rect 104678 382170 104734 382226
rect 104802 382170 104858 382226
rect 104678 382046 104734 382102
rect 104802 382046 104858 382102
rect 104678 381922 104734 381978
rect 104802 381922 104858 381978
rect 135398 382294 135454 382350
rect 135522 382294 135578 382350
rect 135398 382170 135454 382226
rect 135522 382170 135578 382226
rect 135398 382046 135454 382102
rect 135522 382046 135578 382102
rect 135398 381922 135454 381978
rect 135522 381922 135578 381978
rect 166118 382294 166174 382350
rect 166242 382294 166298 382350
rect 166118 382170 166174 382226
rect 166242 382170 166298 382226
rect 166118 382046 166174 382102
rect 166242 382046 166298 382102
rect 166118 381922 166174 381978
rect 166242 381922 166298 381978
rect 196838 382294 196894 382350
rect 196962 382294 197018 382350
rect 196838 382170 196894 382226
rect 196962 382170 197018 382226
rect 196838 382046 196894 382102
rect 196962 382046 197018 382102
rect 196838 381922 196894 381978
rect 196962 381922 197018 381978
rect 227558 382294 227614 382350
rect 227682 382294 227738 382350
rect 227558 382170 227614 382226
rect 227682 382170 227738 382226
rect 227558 382046 227614 382102
rect 227682 382046 227738 382102
rect 227558 381922 227614 381978
rect 227682 381922 227738 381978
rect 258278 382294 258334 382350
rect 258402 382294 258458 382350
rect 258278 382170 258334 382226
rect 258402 382170 258458 382226
rect 258278 382046 258334 382102
rect 258402 382046 258458 382102
rect 258278 381922 258334 381978
rect 258402 381922 258458 381978
rect 288998 382294 289054 382350
rect 289122 382294 289178 382350
rect 288998 382170 289054 382226
rect 289122 382170 289178 382226
rect 288998 382046 289054 382102
rect 289122 382046 289178 382102
rect 288998 381922 289054 381978
rect 289122 381922 289178 381978
rect 319718 382294 319774 382350
rect 319842 382294 319898 382350
rect 319718 382170 319774 382226
rect 319842 382170 319898 382226
rect 319718 382046 319774 382102
rect 319842 382046 319898 382102
rect 319718 381922 319774 381978
rect 319842 381922 319898 381978
rect 350438 382294 350494 382350
rect 350562 382294 350618 382350
rect 350438 382170 350494 382226
rect 350562 382170 350618 382226
rect 350438 382046 350494 382102
rect 350562 382046 350618 382102
rect 350438 381922 350494 381978
rect 350562 381922 350618 381978
rect 381158 382294 381214 382350
rect 381282 382294 381338 382350
rect 381158 382170 381214 382226
rect 381282 382170 381338 382226
rect 381158 382046 381214 382102
rect 381282 382046 381338 382102
rect 381158 381922 381214 381978
rect 381282 381922 381338 381978
rect 411878 382294 411934 382350
rect 412002 382294 412058 382350
rect 411878 382170 411934 382226
rect 412002 382170 412058 382226
rect 411878 382046 411934 382102
rect 412002 382046 412058 382102
rect 411878 381922 411934 381978
rect 412002 381922 412058 381978
rect 442598 382294 442654 382350
rect 442722 382294 442778 382350
rect 442598 382170 442654 382226
rect 442722 382170 442778 382226
rect 442598 382046 442654 382102
rect 442722 382046 442778 382102
rect 442598 381922 442654 381978
rect 442722 381922 442778 381978
rect 473318 382294 473374 382350
rect 473442 382294 473498 382350
rect 473318 382170 473374 382226
rect 473442 382170 473498 382226
rect 473318 382046 473374 382102
rect 473442 382046 473498 382102
rect 473318 381922 473374 381978
rect 473442 381922 473498 381978
rect 504038 382294 504094 382350
rect 504162 382294 504218 382350
rect 504038 382170 504094 382226
rect 504162 382170 504218 382226
rect 504038 382046 504094 382102
rect 504162 382046 504218 382102
rect 504038 381922 504094 381978
rect 504162 381922 504218 381978
rect 534758 382294 534814 382350
rect 534882 382294 534938 382350
rect 534758 382170 534814 382226
rect 534882 382170 534938 382226
rect 534758 382046 534814 382102
rect 534882 382046 534938 382102
rect 534758 381922 534814 381978
rect 534882 381922 534938 381978
rect 565478 382294 565534 382350
rect 565602 382294 565658 382350
rect 565478 382170 565534 382226
rect 565602 382170 565658 382226
rect 565478 382046 565534 382102
rect 565602 382046 565658 382102
rect 565478 381922 565534 381978
rect 565602 381922 565658 381978
rect 5514 364294 5570 364350
rect 5638 364294 5694 364350
rect 5762 364294 5818 364350
rect 5886 364294 5942 364350
rect 5514 364170 5570 364226
rect 5638 364170 5694 364226
rect 5762 364170 5818 364226
rect 5886 364170 5942 364226
rect 5514 364046 5570 364102
rect 5638 364046 5694 364102
rect 5762 364046 5818 364102
rect 5886 364046 5942 364102
rect 5514 363922 5570 363978
rect 5638 363922 5694 363978
rect 5762 363922 5818 363978
rect 5886 363922 5942 363978
rect -860 346294 -804 346350
rect -736 346294 -680 346350
rect -612 346294 -556 346350
rect -488 346294 -432 346350
rect -860 346170 -804 346226
rect -736 346170 -680 346226
rect -612 346170 -556 346226
rect -488 346170 -432 346226
rect -860 346046 -804 346102
rect -736 346046 -680 346102
rect -612 346046 -556 346102
rect -488 346046 -432 346102
rect -860 345922 -804 345978
rect -736 345922 -680 345978
rect -612 345922 -556 345978
rect -488 345922 -432 345978
rect 27878 370294 27934 370350
rect 28002 370294 28058 370350
rect 27878 370170 27934 370226
rect 28002 370170 28058 370226
rect 27878 370046 27934 370102
rect 28002 370046 28058 370102
rect 27878 369922 27934 369978
rect 28002 369922 28058 369978
rect 58598 370294 58654 370350
rect 58722 370294 58778 370350
rect 58598 370170 58654 370226
rect 58722 370170 58778 370226
rect 58598 370046 58654 370102
rect 58722 370046 58778 370102
rect 58598 369922 58654 369978
rect 58722 369922 58778 369978
rect 89318 370294 89374 370350
rect 89442 370294 89498 370350
rect 89318 370170 89374 370226
rect 89442 370170 89498 370226
rect 89318 370046 89374 370102
rect 89442 370046 89498 370102
rect 89318 369922 89374 369978
rect 89442 369922 89498 369978
rect 120038 370294 120094 370350
rect 120162 370294 120218 370350
rect 120038 370170 120094 370226
rect 120162 370170 120218 370226
rect 120038 370046 120094 370102
rect 120162 370046 120218 370102
rect 120038 369922 120094 369978
rect 120162 369922 120218 369978
rect 150758 370294 150814 370350
rect 150882 370294 150938 370350
rect 150758 370170 150814 370226
rect 150882 370170 150938 370226
rect 150758 370046 150814 370102
rect 150882 370046 150938 370102
rect 150758 369922 150814 369978
rect 150882 369922 150938 369978
rect 181478 370294 181534 370350
rect 181602 370294 181658 370350
rect 181478 370170 181534 370226
rect 181602 370170 181658 370226
rect 181478 370046 181534 370102
rect 181602 370046 181658 370102
rect 181478 369922 181534 369978
rect 181602 369922 181658 369978
rect 212198 370294 212254 370350
rect 212322 370294 212378 370350
rect 212198 370170 212254 370226
rect 212322 370170 212378 370226
rect 212198 370046 212254 370102
rect 212322 370046 212378 370102
rect 212198 369922 212254 369978
rect 212322 369922 212378 369978
rect 242918 370294 242974 370350
rect 243042 370294 243098 370350
rect 242918 370170 242974 370226
rect 243042 370170 243098 370226
rect 242918 370046 242974 370102
rect 243042 370046 243098 370102
rect 242918 369922 242974 369978
rect 243042 369922 243098 369978
rect 273638 370294 273694 370350
rect 273762 370294 273818 370350
rect 273638 370170 273694 370226
rect 273762 370170 273818 370226
rect 273638 370046 273694 370102
rect 273762 370046 273818 370102
rect 273638 369922 273694 369978
rect 273762 369922 273818 369978
rect 304358 370294 304414 370350
rect 304482 370294 304538 370350
rect 304358 370170 304414 370226
rect 304482 370170 304538 370226
rect 304358 370046 304414 370102
rect 304482 370046 304538 370102
rect 304358 369922 304414 369978
rect 304482 369922 304538 369978
rect 335078 370294 335134 370350
rect 335202 370294 335258 370350
rect 335078 370170 335134 370226
rect 335202 370170 335258 370226
rect 335078 370046 335134 370102
rect 335202 370046 335258 370102
rect 335078 369922 335134 369978
rect 335202 369922 335258 369978
rect 365798 370294 365854 370350
rect 365922 370294 365978 370350
rect 365798 370170 365854 370226
rect 365922 370170 365978 370226
rect 365798 370046 365854 370102
rect 365922 370046 365978 370102
rect 365798 369922 365854 369978
rect 365922 369922 365978 369978
rect 396518 370294 396574 370350
rect 396642 370294 396698 370350
rect 396518 370170 396574 370226
rect 396642 370170 396698 370226
rect 396518 370046 396574 370102
rect 396642 370046 396698 370102
rect 396518 369922 396574 369978
rect 396642 369922 396698 369978
rect 427238 370294 427294 370350
rect 427362 370294 427418 370350
rect 427238 370170 427294 370226
rect 427362 370170 427418 370226
rect 427238 370046 427294 370102
rect 427362 370046 427418 370102
rect 427238 369922 427294 369978
rect 427362 369922 427418 369978
rect 457958 370294 458014 370350
rect 458082 370294 458138 370350
rect 457958 370170 458014 370226
rect 458082 370170 458138 370226
rect 457958 370046 458014 370102
rect 458082 370046 458138 370102
rect 457958 369922 458014 369978
rect 458082 369922 458138 369978
rect 488678 370294 488734 370350
rect 488802 370294 488858 370350
rect 488678 370170 488734 370226
rect 488802 370170 488858 370226
rect 488678 370046 488734 370102
rect 488802 370046 488858 370102
rect 488678 369922 488734 369978
rect 488802 369922 488858 369978
rect 519398 370294 519454 370350
rect 519522 370294 519578 370350
rect 519398 370170 519454 370226
rect 519522 370170 519578 370226
rect 519398 370046 519454 370102
rect 519522 370046 519578 370102
rect 519398 369922 519454 369978
rect 519522 369922 519578 369978
rect 550118 370294 550174 370350
rect 550242 370294 550298 370350
rect 550118 370170 550174 370226
rect 550242 370170 550298 370226
rect 550118 370046 550174 370102
rect 550242 370046 550298 370102
rect 550118 369922 550174 369978
rect 550242 369922 550298 369978
rect 12518 364294 12574 364350
rect 12642 364294 12698 364350
rect 12518 364170 12574 364226
rect 12642 364170 12698 364226
rect 12518 364046 12574 364102
rect 12642 364046 12698 364102
rect 12518 363922 12574 363978
rect 12642 363922 12698 363978
rect 43238 364294 43294 364350
rect 43362 364294 43418 364350
rect 43238 364170 43294 364226
rect 43362 364170 43418 364226
rect 43238 364046 43294 364102
rect 43362 364046 43418 364102
rect 43238 363922 43294 363978
rect 43362 363922 43418 363978
rect 73958 364294 74014 364350
rect 74082 364294 74138 364350
rect 73958 364170 74014 364226
rect 74082 364170 74138 364226
rect 73958 364046 74014 364102
rect 74082 364046 74138 364102
rect 73958 363922 74014 363978
rect 74082 363922 74138 363978
rect 104678 364294 104734 364350
rect 104802 364294 104858 364350
rect 104678 364170 104734 364226
rect 104802 364170 104858 364226
rect 104678 364046 104734 364102
rect 104802 364046 104858 364102
rect 104678 363922 104734 363978
rect 104802 363922 104858 363978
rect 135398 364294 135454 364350
rect 135522 364294 135578 364350
rect 135398 364170 135454 364226
rect 135522 364170 135578 364226
rect 135398 364046 135454 364102
rect 135522 364046 135578 364102
rect 135398 363922 135454 363978
rect 135522 363922 135578 363978
rect 166118 364294 166174 364350
rect 166242 364294 166298 364350
rect 166118 364170 166174 364226
rect 166242 364170 166298 364226
rect 166118 364046 166174 364102
rect 166242 364046 166298 364102
rect 166118 363922 166174 363978
rect 166242 363922 166298 363978
rect 196838 364294 196894 364350
rect 196962 364294 197018 364350
rect 196838 364170 196894 364226
rect 196962 364170 197018 364226
rect 196838 364046 196894 364102
rect 196962 364046 197018 364102
rect 196838 363922 196894 363978
rect 196962 363922 197018 363978
rect 227558 364294 227614 364350
rect 227682 364294 227738 364350
rect 227558 364170 227614 364226
rect 227682 364170 227738 364226
rect 227558 364046 227614 364102
rect 227682 364046 227738 364102
rect 227558 363922 227614 363978
rect 227682 363922 227738 363978
rect 258278 364294 258334 364350
rect 258402 364294 258458 364350
rect 258278 364170 258334 364226
rect 258402 364170 258458 364226
rect 258278 364046 258334 364102
rect 258402 364046 258458 364102
rect 258278 363922 258334 363978
rect 258402 363922 258458 363978
rect 288998 364294 289054 364350
rect 289122 364294 289178 364350
rect 288998 364170 289054 364226
rect 289122 364170 289178 364226
rect 288998 364046 289054 364102
rect 289122 364046 289178 364102
rect 288998 363922 289054 363978
rect 289122 363922 289178 363978
rect 319718 364294 319774 364350
rect 319842 364294 319898 364350
rect 319718 364170 319774 364226
rect 319842 364170 319898 364226
rect 319718 364046 319774 364102
rect 319842 364046 319898 364102
rect 319718 363922 319774 363978
rect 319842 363922 319898 363978
rect 350438 364294 350494 364350
rect 350562 364294 350618 364350
rect 350438 364170 350494 364226
rect 350562 364170 350618 364226
rect 350438 364046 350494 364102
rect 350562 364046 350618 364102
rect 350438 363922 350494 363978
rect 350562 363922 350618 363978
rect 381158 364294 381214 364350
rect 381282 364294 381338 364350
rect 381158 364170 381214 364226
rect 381282 364170 381338 364226
rect 381158 364046 381214 364102
rect 381282 364046 381338 364102
rect 381158 363922 381214 363978
rect 381282 363922 381338 363978
rect 411878 364294 411934 364350
rect 412002 364294 412058 364350
rect 411878 364170 411934 364226
rect 412002 364170 412058 364226
rect 411878 364046 411934 364102
rect 412002 364046 412058 364102
rect 411878 363922 411934 363978
rect 412002 363922 412058 363978
rect 442598 364294 442654 364350
rect 442722 364294 442778 364350
rect 442598 364170 442654 364226
rect 442722 364170 442778 364226
rect 442598 364046 442654 364102
rect 442722 364046 442778 364102
rect 442598 363922 442654 363978
rect 442722 363922 442778 363978
rect 473318 364294 473374 364350
rect 473442 364294 473498 364350
rect 473318 364170 473374 364226
rect 473442 364170 473498 364226
rect 473318 364046 473374 364102
rect 473442 364046 473498 364102
rect 473318 363922 473374 363978
rect 473442 363922 473498 363978
rect 504038 364294 504094 364350
rect 504162 364294 504218 364350
rect 504038 364170 504094 364226
rect 504162 364170 504218 364226
rect 504038 364046 504094 364102
rect 504162 364046 504218 364102
rect 504038 363922 504094 363978
rect 504162 363922 504218 363978
rect 534758 364294 534814 364350
rect 534882 364294 534938 364350
rect 534758 364170 534814 364226
rect 534882 364170 534938 364226
rect 534758 364046 534814 364102
rect 534882 364046 534938 364102
rect 534758 363922 534814 363978
rect 534882 363922 534938 363978
rect 565478 364294 565534 364350
rect 565602 364294 565658 364350
rect 565478 364170 565534 364226
rect 565602 364170 565658 364226
rect 565478 364046 565534 364102
rect 565602 364046 565658 364102
rect 565478 363922 565534 363978
rect 565602 363922 565658 363978
rect 589194 400294 589250 400350
rect 589318 400294 589374 400350
rect 589442 400294 589498 400350
rect 589566 400294 589622 400350
rect 589194 400170 589250 400226
rect 589318 400170 589374 400226
rect 589442 400170 589498 400226
rect 589566 400170 589622 400226
rect 589194 400046 589250 400102
rect 589318 400046 589374 400102
rect 589442 400046 589498 400102
rect 589566 400046 589622 400102
rect 589194 399922 589250 399978
rect 589318 399922 589374 399978
rect 589442 399922 589498 399978
rect 589566 399922 589622 399978
rect 589194 382294 589250 382350
rect 589318 382294 589374 382350
rect 589442 382294 589498 382350
rect 589566 382294 589622 382350
rect 589194 382170 589250 382226
rect 589318 382170 589374 382226
rect 589442 382170 589498 382226
rect 589566 382170 589622 382226
rect 589194 382046 589250 382102
rect 589318 382046 589374 382102
rect 589442 382046 589498 382102
rect 589566 382046 589622 382102
rect 589194 381922 589250 381978
rect 589318 381922 589374 381978
rect 589442 381922 589498 381978
rect 589566 381922 589622 381978
rect 27878 352294 27934 352350
rect 28002 352294 28058 352350
rect 27878 352170 27934 352226
rect 28002 352170 28058 352226
rect 27878 352046 27934 352102
rect 28002 352046 28058 352102
rect 27878 351922 27934 351978
rect 28002 351922 28058 351978
rect 58598 352294 58654 352350
rect 58722 352294 58778 352350
rect 58598 352170 58654 352226
rect 58722 352170 58778 352226
rect 58598 352046 58654 352102
rect 58722 352046 58778 352102
rect 58598 351922 58654 351978
rect 58722 351922 58778 351978
rect 89318 352294 89374 352350
rect 89442 352294 89498 352350
rect 89318 352170 89374 352226
rect 89442 352170 89498 352226
rect 89318 352046 89374 352102
rect 89442 352046 89498 352102
rect 89318 351922 89374 351978
rect 89442 351922 89498 351978
rect 120038 352294 120094 352350
rect 120162 352294 120218 352350
rect 120038 352170 120094 352226
rect 120162 352170 120218 352226
rect 120038 352046 120094 352102
rect 120162 352046 120218 352102
rect 120038 351922 120094 351978
rect 120162 351922 120218 351978
rect 150758 352294 150814 352350
rect 150882 352294 150938 352350
rect 150758 352170 150814 352226
rect 150882 352170 150938 352226
rect 150758 352046 150814 352102
rect 150882 352046 150938 352102
rect 150758 351922 150814 351978
rect 150882 351922 150938 351978
rect 181478 352294 181534 352350
rect 181602 352294 181658 352350
rect 181478 352170 181534 352226
rect 181602 352170 181658 352226
rect 181478 352046 181534 352102
rect 181602 352046 181658 352102
rect 181478 351922 181534 351978
rect 181602 351922 181658 351978
rect 212198 352294 212254 352350
rect 212322 352294 212378 352350
rect 212198 352170 212254 352226
rect 212322 352170 212378 352226
rect 212198 352046 212254 352102
rect 212322 352046 212378 352102
rect 212198 351922 212254 351978
rect 212322 351922 212378 351978
rect 242918 352294 242974 352350
rect 243042 352294 243098 352350
rect 242918 352170 242974 352226
rect 243042 352170 243098 352226
rect 242918 352046 242974 352102
rect 243042 352046 243098 352102
rect 242918 351922 242974 351978
rect 243042 351922 243098 351978
rect 273638 352294 273694 352350
rect 273762 352294 273818 352350
rect 273638 352170 273694 352226
rect 273762 352170 273818 352226
rect 273638 352046 273694 352102
rect 273762 352046 273818 352102
rect 273638 351922 273694 351978
rect 273762 351922 273818 351978
rect 304358 352294 304414 352350
rect 304482 352294 304538 352350
rect 304358 352170 304414 352226
rect 304482 352170 304538 352226
rect 304358 352046 304414 352102
rect 304482 352046 304538 352102
rect 304358 351922 304414 351978
rect 304482 351922 304538 351978
rect 335078 352294 335134 352350
rect 335202 352294 335258 352350
rect 335078 352170 335134 352226
rect 335202 352170 335258 352226
rect 335078 352046 335134 352102
rect 335202 352046 335258 352102
rect 335078 351922 335134 351978
rect 335202 351922 335258 351978
rect 365798 352294 365854 352350
rect 365922 352294 365978 352350
rect 365798 352170 365854 352226
rect 365922 352170 365978 352226
rect 365798 352046 365854 352102
rect 365922 352046 365978 352102
rect 365798 351922 365854 351978
rect 365922 351922 365978 351978
rect 396518 352294 396574 352350
rect 396642 352294 396698 352350
rect 396518 352170 396574 352226
rect 396642 352170 396698 352226
rect 396518 352046 396574 352102
rect 396642 352046 396698 352102
rect 396518 351922 396574 351978
rect 396642 351922 396698 351978
rect 427238 352294 427294 352350
rect 427362 352294 427418 352350
rect 427238 352170 427294 352226
rect 427362 352170 427418 352226
rect 427238 352046 427294 352102
rect 427362 352046 427418 352102
rect 427238 351922 427294 351978
rect 427362 351922 427418 351978
rect 457958 352294 458014 352350
rect 458082 352294 458138 352350
rect 457958 352170 458014 352226
rect 458082 352170 458138 352226
rect 457958 352046 458014 352102
rect 458082 352046 458138 352102
rect 457958 351922 458014 351978
rect 458082 351922 458138 351978
rect 488678 352294 488734 352350
rect 488802 352294 488858 352350
rect 488678 352170 488734 352226
rect 488802 352170 488858 352226
rect 488678 352046 488734 352102
rect 488802 352046 488858 352102
rect 488678 351922 488734 351978
rect 488802 351922 488858 351978
rect 519398 352294 519454 352350
rect 519522 352294 519578 352350
rect 519398 352170 519454 352226
rect 519522 352170 519578 352226
rect 519398 352046 519454 352102
rect 519522 352046 519578 352102
rect 519398 351922 519454 351978
rect 519522 351922 519578 351978
rect 550118 352294 550174 352350
rect 550242 352294 550298 352350
rect 550118 352170 550174 352226
rect 550242 352170 550298 352226
rect 550118 352046 550174 352102
rect 550242 352046 550298 352102
rect 550118 351922 550174 351978
rect 550242 351922 550298 351978
rect 5514 346294 5570 346350
rect 5638 346294 5694 346350
rect 5762 346294 5818 346350
rect 5886 346294 5942 346350
rect 5514 346170 5570 346226
rect 5638 346170 5694 346226
rect 5762 346170 5818 346226
rect 5886 346170 5942 346226
rect 5514 346046 5570 346102
rect 5638 346046 5694 346102
rect 5762 346046 5818 346102
rect 5886 346046 5942 346102
rect 5514 345922 5570 345978
rect 5638 345922 5694 345978
rect 5762 345922 5818 345978
rect 5886 345922 5942 345978
rect -860 328294 -804 328350
rect -736 328294 -680 328350
rect -612 328294 -556 328350
rect -488 328294 -432 328350
rect -860 328170 -804 328226
rect -736 328170 -680 328226
rect -612 328170 -556 328226
rect -488 328170 -432 328226
rect -860 328046 -804 328102
rect -736 328046 -680 328102
rect -612 328046 -556 328102
rect -488 328046 -432 328102
rect -860 327922 -804 327978
rect -736 327922 -680 327978
rect -612 327922 -556 327978
rect -488 327922 -432 327978
rect 12518 346294 12574 346350
rect 12642 346294 12698 346350
rect 12518 346170 12574 346226
rect 12642 346170 12698 346226
rect 12518 346046 12574 346102
rect 12642 346046 12698 346102
rect 12518 345922 12574 345978
rect 12642 345922 12698 345978
rect 43238 346294 43294 346350
rect 43362 346294 43418 346350
rect 43238 346170 43294 346226
rect 43362 346170 43418 346226
rect 43238 346046 43294 346102
rect 43362 346046 43418 346102
rect 43238 345922 43294 345978
rect 43362 345922 43418 345978
rect 73958 346294 74014 346350
rect 74082 346294 74138 346350
rect 73958 346170 74014 346226
rect 74082 346170 74138 346226
rect 73958 346046 74014 346102
rect 74082 346046 74138 346102
rect 73958 345922 74014 345978
rect 74082 345922 74138 345978
rect 104678 346294 104734 346350
rect 104802 346294 104858 346350
rect 104678 346170 104734 346226
rect 104802 346170 104858 346226
rect 104678 346046 104734 346102
rect 104802 346046 104858 346102
rect 104678 345922 104734 345978
rect 104802 345922 104858 345978
rect 135398 346294 135454 346350
rect 135522 346294 135578 346350
rect 135398 346170 135454 346226
rect 135522 346170 135578 346226
rect 135398 346046 135454 346102
rect 135522 346046 135578 346102
rect 135398 345922 135454 345978
rect 135522 345922 135578 345978
rect 166118 346294 166174 346350
rect 166242 346294 166298 346350
rect 166118 346170 166174 346226
rect 166242 346170 166298 346226
rect 166118 346046 166174 346102
rect 166242 346046 166298 346102
rect 166118 345922 166174 345978
rect 166242 345922 166298 345978
rect 196838 346294 196894 346350
rect 196962 346294 197018 346350
rect 196838 346170 196894 346226
rect 196962 346170 197018 346226
rect 196838 346046 196894 346102
rect 196962 346046 197018 346102
rect 196838 345922 196894 345978
rect 196962 345922 197018 345978
rect 227558 346294 227614 346350
rect 227682 346294 227738 346350
rect 227558 346170 227614 346226
rect 227682 346170 227738 346226
rect 227558 346046 227614 346102
rect 227682 346046 227738 346102
rect 227558 345922 227614 345978
rect 227682 345922 227738 345978
rect 258278 346294 258334 346350
rect 258402 346294 258458 346350
rect 258278 346170 258334 346226
rect 258402 346170 258458 346226
rect 258278 346046 258334 346102
rect 258402 346046 258458 346102
rect 258278 345922 258334 345978
rect 258402 345922 258458 345978
rect 288998 346294 289054 346350
rect 289122 346294 289178 346350
rect 288998 346170 289054 346226
rect 289122 346170 289178 346226
rect 288998 346046 289054 346102
rect 289122 346046 289178 346102
rect 288998 345922 289054 345978
rect 289122 345922 289178 345978
rect 319718 346294 319774 346350
rect 319842 346294 319898 346350
rect 319718 346170 319774 346226
rect 319842 346170 319898 346226
rect 319718 346046 319774 346102
rect 319842 346046 319898 346102
rect 319718 345922 319774 345978
rect 319842 345922 319898 345978
rect 350438 346294 350494 346350
rect 350562 346294 350618 346350
rect 350438 346170 350494 346226
rect 350562 346170 350618 346226
rect 350438 346046 350494 346102
rect 350562 346046 350618 346102
rect 350438 345922 350494 345978
rect 350562 345922 350618 345978
rect 381158 346294 381214 346350
rect 381282 346294 381338 346350
rect 381158 346170 381214 346226
rect 381282 346170 381338 346226
rect 381158 346046 381214 346102
rect 381282 346046 381338 346102
rect 381158 345922 381214 345978
rect 381282 345922 381338 345978
rect 411878 346294 411934 346350
rect 412002 346294 412058 346350
rect 411878 346170 411934 346226
rect 412002 346170 412058 346226
rect 411878 346046 411934 346102
rect 412002 346046 412058 346102
rect 411878 345922 411934 345978
rect 412002 345922 412058 345978
rect 442598 346294 442654 346350
rect 442722 346294 442778 346350
rect 442598 346170 442654 346226
rect 442722 346170 442778 346226
rect 442598 346046 442654 346102
rect 442722 346046 442778 346102
rect 442598 345922 442654 345978
rect 442722 345922 442778 345978
rect 473318 346294 473374 346350
rect 473442 346294 473498 346350
rect 473318 346170 473374 346226
rect 473442 346170 473498 346226
rect 473318 346046 473374 346102
rect 473442 346046 473498 346102
rect 473318 345922 473374 345978
rect 473442 345922 473498 345978
rect 504038 346294 504094 346350
rect 504162 346294 504218 346350
rect 504038 346170 504094 346226
rect 504162 346170 504218 346226
rect 504038 346046 504094 346102
rect 504162 346046 504218 346102
rect 504038 345922 504094 345978
rect 504162 345922 504218 345978
rect 534758 346294 534814 346350
rect 534882 346294 534938 346350
rect 534758 346170 534814 346226
rect 534882 346170 534938 346226
rect 534758 346046 534814 346102
rect 534882 346046 534938 346102
rect 534758 345922 534814 345978
rect 534882 345922 534938 345978
rect 565478 346294 565534 346350
rect 565602 346294 565658 346350
rect 565478 346170 565534 346226
rect 565602 346170 565658 346226
rect 565478 346046 565534 346102
rect 565602 346046 565658 346102
rect 565478 345922 565534 345978
rect 565602 345922 565658 345978
rect 27878 334294 27934 334350
rect 28002 334294 28058 334350
rect 27878 334170 27934 334226
rect 28002 334170 28058 334226
rect 27878 334046 27934 334102
rect 28002 334046 28058 334102
rect 27878 333922 27934 333978
rect 28002 333922 28058 333978
rect 58598 334294 58654 334350
rect 58722 334294 58778 334350
rect 58598 334170 58654 334226
rect 58722 334170 58778 334226
rect 58598 334046 58654 334102
rect 58722 334046 58778 334102
rect 58598 333922 58654 333978
rect 58722 333922 58778 333978
rect 89318 334294 89374 334350
rect 89442 334294 89498 334350
rect 89318 334170 89374 334226
rect 89442 334170 89498 334226
rect 89318 334046 89374 334102
rect 89442 334046 89498 334102
rect 89318 333922 89374 333978
rect 89442 333922 89498 333978
rect 120038 334294 120094 334350
rect 120162 334294 120218 334350
rect 120038 334170 120094 334226
rect 120162 334170 120218 334226
rect 120038 334046 120094 334102
rect 120162 334046 120218 334102
rect 120038 333922 120094 333978
rect 120162 333922 120218 333978
rect 150758 334294 150814 334350
rect 150882 334294 150938 334350
rect 150758 334170 150814 334226
rect 150882 334170 150938 334226
rect 150758 334046 150814 334102
rect 150882 334046 150938 334102
rect 150758 333922 150814 333978
rect 150882 333922 150938 333978
rect 181478 334294 181534 334350
rect 181602 334294 181658 334350
rect 181478 334170 181534 334226
rect 181602 334170 181658 334226
rect 181478 334046 181534 334102
rect 181602 334046 181658 334102
rect 181478 333922 181534 333978
rect 181602 333922 181658 333978
rect 212198 334294 212254 334350
rect 212322 334294 212378 334350
rect 212198 334170 212254 334226
rect 212322 334170 212378 334226
rect 212198 334046 212254 334102
rect 212322 334046 212378 334102
rect 212198 333922 212254 333978
rect 212322 333922 212378 333978
rect 242918 334294 242974 334350
rect 243042 334294 243098 334350
rect 242918 334170 242974 334226
rect 243042 334170 243098 334226
rect 242918 334046 242974 334102
rect 243042 334046 243098 334102
rect 242918 333922 242974 333978
rect 243042 333922 243098 333978
rect 273638 334294 273694 334350
rect 273762 334294 273818 334350
rect 273638 334170 273694 334226
rect 273762 334170 273818 334226
rect 273638 334046 273694 334102
rect 273762 334046 273818 334102
rect 273638 333922 273694 333978
rect 273762 333922 273818 333978
rect 304358 334294 304414 334350
rect 304482 334294 304538 334350
rect 304358 334170 304414 334226
rect 304482 334170 304538 334226
rect 304358 334046 304414 334102
rect 304482 334046 304538 334102
rect 304358 333922 304414 333978
rect 304482 333922 304538 333978
rect 335078 334294 335134 334350
rect 335202 334294 335258 334350
rect 335078 334170 335134 334226
rect 335202 334170 335258 334226
rect 335078 334046 335134 334102
rect 335202 334046 335258 334102
rect 335078 333922 335134 333978
rect 335202 333922 335258 333978
rect 365798 334294 365854 334350
rect 365922 334294 365978 334350
rect 365798 334170 365854 334226
rect 365922 334170 365978 334226
rect 365798 334046 365854 334102
rect 365922 334046 365978 334102
rect 365798 333922 365854 333978
rect 365922 333922 365978 333978
rect 396518 334294 396574 334350
rect 396642 334294 396698 334350
rect 396518 334170 396574 334226
rect 396642 334170 396698 334226
rect 396518 334046 396574 334102
rect 396642 334046 396698 334102
rect 396518 333922 396574 333978
rect 396642 333922 396698 333978
rect 427238 334294 427294 334350
rect 427362 334294 427418 334350
rect 427238 334170 427294 334226
rect 427362 334170 427418 334226
rect 427238 334046 427294 334102
rect 427362 334046 427418 334102
rect 427238 333922 427294 333978
rect 427362 333922 427418 333978
rect 457958 334294 458014 334350
rect 458082 334294 458138 334350
rect 457958 334170 458014 334226
rect 458082 334170 458138 334226
rect 457958 334046 458014 334102
rect 458082 334046 458138 334102
rect 457958 333922 458014 333978
rect 458082 333922 458138 333978
rect 488678 334294 488734 334350
rect 488802 334294 488858 334350
rect 488678 334170 488734 334226
rect 488802 334170 488858 334226
rect 488678 334046 488734 334102
rect 488802 334046 488858 334102
rect 488678 333922 488734 333978
rect 488802 333922 488858 333978
rect 519398 334294 519454 334350
rect 519522 334294 519578 334350
rect 519398 334170 519454 334226
rect 519522 334170 519578 334226
rect 519398 334046 519454 334102
rect 519522 334046 519578 334102
rect 519398 333922 519454 333978
rect 519522 333922 519578 333978
rect 550118 334294 550174 334350
rect 550242 334294 550298 334350
rect 550118 334170 550174 334226
rect 550242 334170 550298 334226
rect 550118 334046 550174 334102
rect 550242 334046 550298 334102
rect 550118 333922 550174 333978
rect 550242 333922 550298 333978
rect 5514 328294 5570 328350
rect 5638 328294 5694 328350
rect 5762 328294 5818 328350
rect 5886 328294 5942 328350
rect 5514 328170 5570 328226
rect 5638 328170 5694 328226
rect 5762 328170 5818 328226
rect 5886 328170 5942 328226
rect 5514 328046 5570 328102
rect 5638 328046 5694 328102
rect 5762 328046 5818 328102
rect 5886 328046 5942 328102
rect 5514 327922 5570 327978
rect 5638 327922 5694 327978
rect 5762 327922 5818 327978
rect 5886 327922 5942 327978
rect -860 310294 -804 310350
rect -736 310294 -680 310350
rect -612 310294 -556 310350
rect -488 310294 -432 310350
rect -860 310170 -804 310226
rect -736 310170 -680 310226
rect -612 310170 -556 310226
rect -488 310170 -432 310226
rect -860 310046 -804 310102
rect -736 310046 -680 310102
rect -612 310046 -556 310102
rect -488 310046 -432 310102
rect -860 309922 -804 309978
rect -736 309922 -680 309978
rect -612 309922 -556 309978
rect -488 309922 -432 309978
rect 12518 328294 12574 328350
rect 12642 328294 12698 328350
rect 12518 328170 12574 328226
rect 12642 328170 12698 328226
rect 12518 328046 12574 328102
rect 12642 328046 12698 328102
rect 12518 327922 12574 327978
rect 12642 327922 12698 327978
rect 43238 328294 43294 328350
rect 43362 328294 43418 328350
rect 43238 328170 43294 328226
rect 43362 328170 43418 328226
rect 43238 328046 43294 328102
rect 43362 328046 43418 328102
rect 43238 327922 43294 327978
rect 43362 327922 43418 327978
rect 73958 328294 74014 328350
rect 74082 328294 74138 328350
rect 73958 328170 74014 328226
rect 74082 328170 74138 328226
rect 73958 328046 74014 328102
rect 74082 328046 74138 328102
rect 73958 327922 74014 327978
rect 74082 327922 74138 327978
rect 104678 328294 104734 328350
rect 104802 328294 104858 328350
rect 104678 328170 104734 328226
rect 104802 328170 104858 328226
rect 104678 328046 104734 328102
rect 104802 328046 104858 328102
rect 104678 327922 104734 327978
rect 104802 327922 104858 327978
rect 135398 328294 135454 328350
rect 135522 328294 135578 328350
rect 135398 328170 135454 328226
rect 135522 328170 135578 328226
rect 135398 328046 135454 328102
rect 135522 328046 135578 328102
rect 135398 327922 135454 327978
rect 135522 327922 135578 327978
rect 166118 328294 166174 328350
rect 166242 328294 166298 328350
rect 166118 328170 166174 328226
rect 166242 328170 166298 328226
rect 166118 328046 166174 328102
rect 166242 328046 166298 328102
rect 166118 327922 166174 327978
rect 166242 327922 166298 327978
rect 196838 328294 196894 328350
rect 196962 328294 197018 328350
rect 196838 328170 196894 328226
rect 196962 328170 197018 328226
rect 196838 328046 196894 328102
rect 196962 328046 197018 328102
rect 196838 327922 196894 327978
rect 196962 327922 197018 327978
rect 227558 328294 227614 328350
rect 227682 328294 227738 328350
rect 227558 328170 227614 328226
rect 227682 328170 227738 328226
rect 227558 328046 227614 328102
rect 227682 328046 227738 328102
rect 227558 327922 227614 327978
rect 227682 327922 227738 327978
rect 258278 328294 258334 328350
rect 258402 328294 258458 328350
rect 258278 328170 258334 328226
rect 258402 328170 258458 328226
rect 258278 328046 258334 328102
rect 258402 328046 258458 328102
rect 258278 327922 258334 327978
rect 258402 327922 258458 327978
rect 288998 328294 289054 328350
rect 289122 328294 289178 328350
rect 288998 328170 289054 328226
rect 289122 328170 289178 328226
rect 288998 328046 289054 328102
rect 289122 328046 289178 328102
rect 288998 327922 289054 327978
rect 289122 327922 289178 327978
rect 319718 328294 319774 328350
rect 319842 328294 319898 328350
rect 319718 328170 319774 328226
rect 319842 328170 319898 328226
rect 319718 328046 319774 328102
rect 319842 328046 319898 328102
rect 319718 327922 319774 327978
rect 319842 327922 319898 327978
rect 350438 328294 350494 328350
rect 350562 328294 350618 328350
rect 350438 328170 350494 328226
rect 350562 328170 350618 328226
rect 350438 328046 350494 328102
rect 350562 328046 350618 328102
rect 350438 327922 350494 327978
rect 350562 327922 350618 327978
rect 381158 328294 381214 328350
rect 381282 328294 381338 328350
rect 381158 328170 381214 328226
rect 381282 328170 381338 328226
rect 381158 328046 381214 328102
rect 381282 328046 381338 328102
rect 381158 327922 381214 327978
rect 381282 327922 381338 327978
rect 411878 328294 411934 328350
rect 412002 328294 412058 328350
rect 411878 328170 411934 328226
rect 412002 328170 412058 328226
rect 411878 328046 411934 328102
rect 412002 328046 412058 328102
rect 411878 327922 411934 327978
rect 412002 327922 412058 327978
rect 442598 328294 442654 328350
rect 442722 328294 442778 328350
rect 442598 328170 442654 328226
rect 442722 328170 442778 328226
rect 442598 328046 442654 328102
rect 442722 328046 442778 328102
rect 442598 327922 442654 327978
rect 442722 327922 442778 327978
rect 473318 328294 473374 328350
rect 473442 328294 473498 328350
rect 473318 328170 473374 328226
rect 473442 328170 473498 328226
rect 473318 328046 473374 328102
rect 473442 328046 473498 328102
rect 473318 327922 473374 327978
rect 473442 327922 473498 327978
rect 504038 328294 504094 328350
rect 504162 328294 504218 328350
rect 504038 328170 504094 328226
rect 504162 328170 504218 328226
rect 504038 328046 504094 328102
rect 504162 328046 504218 328102
rect 504038 327922 504094 327978
rect 504162 327922 504218 327978
rect 534758 328294 534814 328350
rect 534882 328294 534938 328350
rect 534758 328170 534814 328226
rect 534882 328170 534938 328226
rect 534758 328046 534814 328102
rect 534882 328046 534938 328102
rect 534758 327922 534814 327978
rect 534882 327922 534938 327978
rect 565478 328294 565534 328350
rect 565602 328294 565658 328350
rect 565478 328170 565534 328226
rect 565602 328170 565658 328226
rect 565478 328046 565534 328102
rect 565602 328046 565658 328102
rect 565478 327922 565534 327978
rect 565602 327922 565658 327978
rect 589194 364294 589250 364350
rect 589318 364294 589374 364350
rect 589442 364294 589498 364350
rect 589566 364294 589622 364350
rect 589194 364170 589250 364226
rect 589318 364170 589374 364226
rect 589442 364170 589498 364226
rect 589566 364170 589622 364226
rect 589194 364046 589250 364102
rect 589318 364046 589374 364102
rect 589442 364046 589498 364102
rect 589566 364046 589622 364102
rect 592914 424294 592970 424350
rect 593038 424294 593094 424350
rect 593162 424294 593218 424350
rect 593286 424294 593342 424350
rect 592914 424170 592970 424226
rect 593038 424170 593094 424226
rect 593162 424170 593218 424226
rect 593286 424170 593342 424226
rect 592914 424046 592970 424102
rect 593038 424046 593094 424102
rect 593162 424046 593218 424102
rect 593286 424046 593342 424102
rect 592914 423922 592970 423978
rect 593038 423922 593094 423978
rect 593162 423922 593218 423978
rect 593286 423922 593342 423978
rect 592914 406294 592970 406350
rect 593038 406294 593094 406350
rect 593162 406294 593218 406350
rect 593286 406294 593342 406350
rect 592914 406170 592970 406226
rect 593038 406170 593094 406226
rect 593162 406170 593218 406226
rect 593286 406170 593342 406226
rect 592914 406046 592970 406102
rect 593038 406046 593094 406102
rect 593162 406046 593218 406102
rect 593286 406046 593342 406102
rect 592914 405922 592970 405978
rect 593038 405922 593094 405978
rect 593162 405922 593218 405978
rect 593286 405922 593342 405978
rect 592914 388294 592970 388350
rect 593038 388294 593094 388350
rect 593162 388294 593218 388350
rect 593286 388294 593342 388350
rect 592914 388170 592970 388226
rect 593038 388170 593094 388226
rect 593162 388170 593218 388226
rect 593286 388170 593342 388226
rect 592914 388046 592970 388102
rect 593038 388046 593094 388102
rect 593162 388046 593218 388102
rect 593286 388046 593342 388102
rect 592914 387922 592970 387978
rect 593038 387922 593094 387978
rect 593162 387922 593218 387978
rect 593286 387922 593342 387978
rect 592914 370294 592970 370350
rect 593038 370294 593094 370350
rect 593162 370294 593218 370350
rect 593286 370294 593342 370350
rect 592914 370170 592970 370226
rect 593038 370170 593094 370226
rect 593162 370170 593218 370226
rect 593286 370170 593342 370226
rect 592914 370046 592970 370102
rect 593038 370046 593094 370102
rect 593162 370046 593218 370102
rect 593286 370046 593342 370102
rect 592914 369922 592970 369978
rect 593038 369922 593094 369978
rect 593162 369922 593218 369978
rect 593286 369922 593342 369978
rect 589194 363922 589250 363978
rect 589318 363922 589374 363978
rect 589442 363922 589498 363978
rect 589566 363922 589622 363978
rect 589194 346294 589250 346350
rect 589318 346294 589374 346350
rect 589442 346294 589498 346350
rect 589566 346294 589622 346350
rect 589194 346170 589250 346226
rect 589318 346170 589374 346226
rect 589442 346170 589498 346226
rect 589566 346170 589622 346226
rect 589194 346046 589250 346102
rect 589318 346046 589374 346102
rect 589442 346046 589498 346102
rect 589566 346046 589622 346102
rect 589194 345922 589250 345978
rect 589318 345922 589374 345978
rect 589442 345922 589498 345978
rect 589566 345922 589622 345978
rect 27878 316294 27934 316350
rect 28002 316294 28058 316350
rect 27878 316170 27934 316226
rect 28002 316170 28058 316226
rect 27878 316046 27934 316102
rect 28002 316046 28058 316102
rect 27878 315922 27934 315978
rect 28002 315922 28058 315978
rect 58598 316294 58654 316350
rect 58722 316294 58778 316350
rect 58598 316170 58654 316226
rect 58722 316170 58778 316226
rect 58598 316046 58654 316102
rect 58722 316046 58778 316102
rect 58598 315922 58654 315978
rect 58722 315922 58778 315978
rect 89318 316294 89374 316350
rect 89442 316294 89498 316350
rect 89318 316170 89374 316226
rect 89442 316170 89498 316226
rect 89318 316046 89374 316102
rect 89442 316046 89498 316102
rect 89318 315922 89374 315978
rect 89442 315922 89498 315978
rect 120038 316294 120094 316350
rect 120162 316294 120218 316350
rect 120038 316170 120094 316226
rect 120162 316170 120218 316226
rect 120038 316046 120094 316102
rect 120162 316046 120218 316102
rect 120038 315922 120094 315978
rect 120162 315922 120218 315978
rect 150758 316294 150814 316350
rect 150882 316294 150938 316350
rect 150758 316170 150814 316226
rect 150882 316170 150938 316226
rect 150758 316046 150814 316102
rect 150882 316046 150938 316102
rect 150758 315922 150814 315978
rect 150882 315922 150938 315978
rect 181478 316294 181534 316350
rect 181602 316294 181658 316350
rect 181478 316170 181534 316226
rect 181602 316170 181658 316226
rect 181478 316046 181534 316102
rect 181602 316046 181658 316102
rect 181478 315922 181534 315978
rect 181602 315922 181658 315978
rect 212198 316294 212254 316350
rect 212322 316294 212378 316350
rect 212198 316170 212254 316226
rect 212322 316170 212378 316226
rect 212198 316046 212254 316102
rect 212322 316046 212378 316102
rect 212198 315922 212254 315978
rect 212322 315922 212378 315978
rect 242918 316294 242974 316350
rect 243042 316294 243098 316350
rect 242918 316170 242974 316226
rect 243042 316170 243098 316226
rect 242918 316046 242974 316102
rect 243042 316046 243098 316102
rect 242918 315922 242974 315978
rect 243042 315922 243098 315978
rect 273638 316294 273694 316350
rect 273762 316294 273818 316350
rect 273638 316170 273694 316226
rect 273762 316170 273818 316226
rect 273638 316046 273694 316102
rect 273762 316046 273818 316102
rect 273638 315922 273694 315978
rect 273762 315922 273818 315978
rect 304358 316294 304414 316350
rect 304482 316294 304538 316350
rect 304358 316170 304414 316226
rect 304482 316170 304538 316226
rect 304358 316046 304414 316102
rect 304482 316046 304538 316102
rect 304358 315922 304414 315978
rect 304482 315922 304538 315978
rect 335078 316294 335134 316350
rect 335202 316294 335258 316350
rect 335078 316170 335134 316226
rect 335202 316170 335258 316226
rect 335078 316046 335134 316102
rect 335202 316046 335258 316102
rect 335078 315922 335134 315978
rect 335202 315922 335258 315978
rect 365798 316294 365854 316350
rect 365922 316294 365978 316350
rect 365798 316170 365854 316226
rect 365922 316170 365978 316226
rect 365798 316046 365854 316102
rect 365922 316046 365978 316102
rect 365798 315922 365854 315978
rect 365922 315922 365978 315978
rect 396518 316294 396574 316350
rect 396642 316294 396698 316350
rect 396518 316170 396574 316226
rect 396642 316170 396698 316226
rect 396518 316046 396574 316102
rect 396642 316046 396698 316102
rect 396518 315922 396574 315978
rect 396642 315922 396698 315978
rect 427238 316294 427294 316350
rect 427362 316294 427418 316350
rect 427238 316170 427294 316226
rect 427362 316170 427418 316226
rect 427238 316046 427294 316102
rect 427362 316046 427418 316102
rect 427238 315922 427294 315978
rect 427362 315922 427418 315978
rect 457958 316294 458014 316350
rect 458082 316294 458138 316350
rect 457958 316170 458014 316226
rect 458082 316170 458138 316226
rect 457958 316046 458014 316102
rect 458082 316046 458138 316102
rect 457958 315922 458014 315978
rect 458082 315922 458138 315978
rect 488678 316294 488734 316350
rect 488802 316294 488858 316350
rect 488678 316170 488734 316226
rect 488802 316170 488858 316226
rect 488678 316046 488734 316102
rect 488802 316046 488858 316102
rect 488678 315922 488734 315978
rect 488802 315922 488858 315978
rect 519398 316294 519454 316350
rect 519522 316294 519578 316350
rect 519398 316170 519454 316226
rect 519522 316170 519578 316226
rect 519398 316046 519454 316102
rect 519522 316046 519578 316102
rect 519398 315922 519454 315978
rect 519522 315922 519578 315978
rect 550118 316294 550174 316350
rect 550242 316294 550298 316350
rect 550118 316170 550174 316226
rect 550242 316170 550298 316226
rect 550118 316046 550174 316102
rect 550242 316046 550298 316102
rect 550118 315922 550174 315978
rect 550242 315922 550298 315978
rect 5514 310294 5570 310350
rect 5638 310294 5694 310350
rect 5762 310294 5818 310350
rect 5886 310294 5942 310350
rect 5514 310170 5570 310226
rect 5638 310170 5694 310226
rect 5762 310170 5818 310226
rect 5886 310170 5942 310226
rect 5514 310046 5570 310102
rect 5638 310046 5694 310102
rect 5762 310046 5818 310102
rect 5886 310046 5942 310102
rect 5514 309922 5570 309978
rect 5638 309922 5694 309978
rect 5762 309922 5818 309978
rect 5886 309922 5942 309978
rect -860 292294 -804 292350
rect -736 292294 -680 292350
rect -612 292294 -556 292350
rect -488 292294 -432 292350
rect -860 292170 -804 292226
rect -736 292170 -680 292226
rect -612 292170 -556 292226
rect -488 292170 -432 292226
rect -860 292046 -804 292102
rect -736 292046 -680 292102
rect -612 292046 -556 292102
rect -488 292046 -432 292102
rect -860 291922 -804 291978
rect -736 291922 -680 291978
rect -612 291922 -556 291978
rect -488 291922 -432 291978
rect 12518 310294 12574 310350
rect 12642 310294 12698 310350
rect 12518 310170 12574 310226
rect 12642 310170 12698 310226
rect 12518 310046 12574 310102
rect 12642 310046 12698 310102
rect 12518 309922 12574 309978
rect 12642 309922 12698 309978
rect 43238 310294 43294 310350
rect 43362 310294 43418 310350
rect 43238 310170 43294 310226
rect 43362 310170 43418 310226
rect 43238 310046 43294 310102
rect 43362 310046 43418 310102
rect 43238 309922 43294 309978
rect 43362 309922 43418 309978
rect 73958 310294 74014 310350
rect 74082 310294 74138 310350
rect 73958 310170 74014 310226
rect 74082 310170 74138 310226
rect 73958 310046 74014 310102
rect 74082 310046 74138 310102
rect 73958 309922 74014 309978
rect 74082 309922 74138 309978
rect 104678 310294 104734 310350
rect 104802 310294 104858 310350
rect 104678 310170 104734 310226
rect 104802 310170 104858 310226
rect 104678 310046 104734 310102
rect 104802 310046 104858 310102
rect 104678 309922 104734 309978
rect 104802 309922 104858 309978
rect 135398 310294 135454 310350
rect 135522 310294 135578 310350
rect 135398 310170 135454 310226
rect 135522 310170 135578 310226
rect 135398 310046 135454 310102
rect 135522 310046 135578 310102
rect 135398 309922 135454 309978
rect 135522 309922 135578 309978
rect 166118 310294 166174 310350
rect 166242 310294 166298 310350
rect 166118 310170 166174 310226
rect 166242 310170 166298 310226
rect 166118 310046 166174 310102
rect 166242 310046 166298 310102
rect 166118 309922 166174 309978
rect 166242 309922 166298 309978
rect 196838 310294 196894 310350
rect 196962 310294 197018 310350
rect 196838 310170 196894 310226
rect 196962 310170 197018 310226
rect 196838 310046 196894 310102
rect 196962 310046 197018 310102
rect 196838 309922 196894 309978
rect 196962 309922 197018 309978
rect 227558 310294 227614 310350
rect 227682 310294 227738 310350
rect 227558 310170 227614 310226
rect 227682 310170 227738 310226
rect 227558 310046 227614 310102
rect 227682 310046 227738 310102
rect 227558 309922 227614 309978
rect 227682 309922 227738 309978
rect 258278 310294 258334 310350
rect 258402 310294 258458 310350
rect 258278 310170 258334 310226
rect 258402 310170 258458 310226
rect 258278 310046 258334 310102
rect 258402 310046 258458 310102
rect 258278 309922 258334 309978
rect 258402 309922 258458 309978
rect 288998 310294 289054 310350
rect 289122 310294 289178 310350
rect 288998 310170 289054 310226
rect 289122 310170 289178 310226
rect 288998 310046 289054 310102
rect 289122 310046 289178 310102
rect 288998 309922 289054 309978
rect 289122 309922 289178 309978
rect 319718 310294 319774 310350
rect 319842 310294 319898 310350
rect 319718 310170 319774 310226
rect 319842 310170 319898 310226
rect 319718 310046 319774 310102
rect 319842 310046 319898 310102
rect 319718 309922 319774 309978
rect 319842 309922 319898 309978
rect 350438 310294 350494 310350
rect 350562 310294 350618 310350
rect 350438 310170 350494 310226
rect 350562 310170 350618 310226
rect 350438 310046 350494 310102
rect 350562 310046 350618 310102
rect 350438 309922 350494 309978
rect 350562 309922 350618 309978
rect 381158 310294 381214 310350
rect 381282 310294 381338 310350
rect 381158 310170 381214 310226
rect 381282 310170 381338 310226
rect 381158 310046 381214 310102
rect 381282 310046 381338 310102
rect 381158 309922 381214 309978
rect 381282 309922 381338 309978
rect 411878 310294 411934 310350
rect 412002 310294 412058 310350
rect 411878 310170 411934 310226
rect 412002 310170 412058 310226
rect 411878 310046 411934 310102
rect 412002 310046 412058 310102
rect 411878 309922 411934 309978
rect 412002 309922 412058 309978
rect 442598 310294 442654 310350
rect 442722 310294 442778 310350
rect 442598 310170 442654 310226
rect 442722 310170 442778 310226
rect 442598 310046 442654 310102
rect 442722 310046 442778 310102
rect 442598 309922 442654 309978
rect 442722 309922 442778 309978
rect 473318 310294 473374 310350
rect 473442 310294 473498 310350
rect 473318 310170 473374 310226
rect 473442 310170 473498 310226
rect 473318 310046 473374 310102
rect 473442 310046 473498 310102
rect 473318 309922 473374 309978
rect 473442 309922 473498 309978
rect 504038 310294 504094 310350
rect 504162 310294 504218 310350
rect 504038 310170 504094 310226
rect 504162 310170 504218 310226
rect 504038 310046 504094 310102
rect 504162 310046 504218 310102
rect 504038 309922 504094 309978
rect 504162 309922 504218 309978
rect 534758 310294 534814 310350
rect 534882 310294 534938 310350
rect 534758 310170 534814 310226
rect 534882 310170 534938 310226
rect 534758 310046 534814 310102
rect 534882 310046 534938 310102
rect 534758 309922 534814 309978
rect 534882 309922 534938 309978
rect 565478 310294 565534 310350
rect 565602 310294 565658 310350
rect 565478 310170 565534 310226
rect 565602 310170 565658 310226
rect 565478 310046 565534 310102
rect 565602 310046 565658 310102
rect 565478 309922 565534 309978
rect 565602 309922 565658 309978
rect 5514 292294 5570 292350
rect 5638 292294 5694 292350
rect 5762 292294 5818 292350
rect 5886 292294 5942 292350
rect 5514 292170 5570 292226
rect 5638 292170 5694 292226
rect 5762 292170 5818 292226
rect 5886 292170 5942 292226
rect 5514 292046 5570 292102
rect 5638 292046 5694 292102
rect 5762 292046 5818 292102
rect 5886 292046 5942 292102
rect 5514 291922 5570 291978
rect 5638 291922 5694 291978
rect 5762 291922 5818 291978
rect 5886 291922 5942 291978
rect -860 274294 -804 274350
rect -736 274294 -680 274350
rect -612 274294 -556 274350
rect -488 274294 -432 274350
rect -860 274170 -804 274226
rect -736 274170 -680 274226
rect -612 274170 -556 274226
rect -488 274170 -432 274226
rect -860 274046 -804 274102
rect -736 274046 -680 274102
rect -612 274046 -556 274102
rect -488 274046 -432 274102
rect -860 273922 -804 273978
rect -736 273922 -680 273978
rect -612 273922 -556 273978
rect -488 273922 -432 273978
rect 27878 298294 27934 298350
rect 28002 298294 28058 298350
rect 27878 298170 27934 298226
rect 28002 298170 28058 298226
rect 27878 298046 27934 298102
rect 28002 298046 28058 298102
rect 27878 297922 27934 297978
rect 28002 297922 28058 297978
rect 58598 298294 58654 298350
rect 58722 298294 58778 298350
rect 58598 298170 58654 298226
rect 58722 298170 58778 298226
rect 58598 298046 58654 298102
rect 58722 298046 58778 298102
rect 58598 297922 58654 297978
rect 58722 297922 58778 297978
rect 89318 298294 89374 298350
rect 89442 298294 89498 298350
rect 89318 298170 89374 298226
rect 89442 298170 89498 298226
rect 89318 298046 89374 298102
rect 89442 298046 89498 298102
rect 89318 297922 89374 297978
rect 89442 297922 89498 297978
rect 120038 298294 120094 298350
rect 120162 298294 120218 298350
rect 120038 298170 120094 298226
rect 120162 298170 120218 298226
rect 120038 298046 120094 298102
rect 120162 298046 120218 298102
rect 120038 297922 120094 297978
rect 120162 297922 120218 297978
rect 150758 298294 150814 298350
rect 150882 298294 150938 298350
rect 150758 298170 150814 298226
rect 150882 298170 150938 298226
rect 150758 298046 150814 298102
rect 150882 298046 150938 298102
rect 150758 297922 150814 297978
rect 150882 297922 150938 297978
rect 181478 298294 181534 298350
rect 181602 298294 181658 298350
rect 181478 298170 181534 298226
rect 181602 298170 181658 298226
rect 181478 298046 181534 298102
rect 181602 298046 181658 298102
rect 181478 297922 181534 297978
rect 181602 297922 181658 297978
rect 212198 298294 212254 298350
rect 212322 298294 212378 298350
rect 212198 298170 212254 298226
rect 212322 298170 212378 298226
rect 212198 298046 212254 298102
rect 212322 298046 212378 298102
rect 212198 297922 212254 297978
rect 212322 297922 212378 297978
rect 242918 298294 242974 298350
rect 243042 298294 243098 298350
rect 242918 298170 242974 298226
rect 243042 298170 243098 298226
rect 242918 298046 242974 298102
rect 243042 298046 243098 298102
rect 242918 297922 242974 297978
rect 243042 297922 243098 297978
rect 273638 298294 273694 298350
rect 273762 298294 273818 298350
rect 273638 298170 273694 298226
rect 273762 298170 273818 298226
rect 273638 298046 273694 298102
rect 273762 298046 273818 298102
rect 273638 297922 273694 297978
rect 273762 297922 273818 297978
rect 304358 298294 304414 298350
rect 304482 298294 304538 298350
rect 304358 298170 304414 298226
rect 304482 298170 304538 298226
rect 304358 298046 304414 298102
rect 304482 298046 304538 298102
rect 304358 297922 304414 297978
rect 304482 297922 304538 297978
rect 335078 298294 335134 298350
rect 335202 298294 335258 298350
rect 335078 298170 335134 298226
rect 335202 298170 335258 298226
rect 335078 298046 335134 298102
rect 335202 298046 335258 298102
rect 335078 297922 335134 297978
rect 335202 297922 335258 297978
rect 365798 298294 365854 298350
rect 365922 298294 365978 298350
rect 365798 298170 365854 298226
rect 365922 298170 365978 298226
rect 365798 298046 365854 298102
rect 365922 298046 365978 298102
rect 365798 297922 365854 297978
rect 365922 297922 365978 297978
rect 396518 298294 396574 298350
rect 396642 298294 396698 298350
rect 396518 298170 396574 298226
rect 396642 298170 396698 298226
rect 396518 298046 396574 298102
rect 396642 298046 396698 298102
rect 396518 297922 396574 297978
rect 396642 297922 396698 297978
rect 427238 298294 427294 298350
rect 427362 298294 427418 298350
rect 427238 298170 427294 298226
rect 427362 298170 427418 298226
rect 427238 298046 427294 298102
rect 427362 298046 427418 298102
rect 427238 297922 427294 297978
rect 427362 297922 427418 297978
rect 457958 298294 458014 298350
rect 458082 298294 458138 298350
rect 457958 298170 458014 298226
rect 458082 298170 458138 298226
rect 457958 298046 458014 298102
rect 458082 298046 458138 298102
rect 457958 297922 458014 297978
rect 458082 297922 458138 297978
rect 488678 298294 488734 298350
rect 488802 298294 488858 298350
rect 488678 298170 488734 298226
rect 488802 298170 488858 298226
rect 488678 298046 488734 298102
rect 488802 298046 488858 298102
rect 488678 297922 488734 297978
rect 488802 297922 488858 297978
rect 519398 298294 519454 298350
rect 519522 298294 519578 298350
rect 519398 298170 519454 298226
rect 519522 298170 519578 298226
rect 519398 298046 519454 298102
rect 519522 298046 519578 298102
rect 519398 297922 519454 297978
rect 519522 297922 519578 297978
rect 550118 298294 550174 298350
rect 550242 298294 550298 298350
rect 550118 298170 550174 298226
rect 550242 298170 550298 298226
rect 550118 298046 550174 298102
rect 550242 298046 550298 298102
rect 550118 297922 550174 297978
rect 550242 297922 550298 297978
rect 12518 292294 12574 292350
rect 12642 292294 12698 292350
rect 12518 292170 12574 292226
rect 12642 292170 12698 292226
rect 12518 292046 12574 292102
rect 12642 292046 12698 292102
rect 12518 291922 12574 291978
rect 12642 291922 12698 291978
rect 43238 292294 43294 292350
rect 43362 292294 43418 292350
rect 43238 292170 43294 292226
rect 43362 292170 43418 292226
rect 43238 292046 43294 292102
rect 43362 292046 43418 292102
rect 43238 291922 43294 291978
rect 43362 291922 43418 291978
rect 73958 292294 74014 292350
rect 74082 292294 74138 292350
rect 73958 292170 74014 292226
rect 74082 292170 74138 292226
rect 73958 292046 74014 292102
rect 74082 292046 74138 292102
rect 73958 291922 74014 291978
rect 74082 291922 74138 291978
rect 104678 292294 104734 292350
rect 104802 292294 104858 292350
rect 104678 292170 104734 292226
rect 104802 292170 104858 292226
rect 104678 292046 104734 292102
rect 104802 292046 104858 292102
rect 104678 291922 104734 291978
rect 104802 291922 104858 291978
rect 135398 292294 135454 292350
rect 135522 292294 135578 292350
rect 135398 292170 135454 292226
rect 135522 292170 135578 292226
rect 135398 292046 135454 292102
rect 135522 292046 135578 292102
rect 135398 291922 135454 291978
rect 135522 291922 135578 291978
rect 166118 292294 166174 292350
rect 166242 292294 166298 292350
rect 166118 292170 166174 292226
rect 166242 292170 166298 292226
rect 166118 292046 166174 292102
rect 166242 292046 166298 292102
rect 166118 291922 166174 291978
rect 166242 291922 166298 291978
rect 196838 292294 196894 292350
rect 196962 292294 197018 292350
rect 196838 292170 196894 292226
rect 196962 292170 197018 292226
rect 196838 292046 196894 292102
rect 196962 292046 197018 292102
rect 196838 291922 196894 291978
rect 196962 291922 197018 291978
rect 227558 292294 227614 292350
rect 227682 292294 227738 292350
rect 227558 292170 227614 292226
rect 227682 292170 227738 292226
rect 227558 292046 227614 292102
rect 227682 292046 227738 292102
rect 227558 291922 227614 291978
rect 227682 291922 227738 291978
rect 258278 292294 258334 292350
rect 258402 292294 258458 292350
rect 258278 292170 258334 292226
rect 258402 292170 258458 292226
rect 258278 292046 258334 292102
rect 258402 292046 258458 292102
rect 258278 291922 258334 291978
rect 258402 291922 258458 291978
rect 288998 292294 289054 292350
rect 289122 292294 289178 292350
rect 288998 292170 289054 292226
rect 289122 292170 289178 292226
rect 288998 292046 289054 292102
rect 289122 292046 289178 292102
rect 288998 291922 289054 291978
rect 289122 291922 289178 291978
rect 319718 292294 319774 292350
rect 319842 292294 319898 292350
rect 319718 292170 319774 292226
rect 319842 292170 319898 292226
rect 319718 292046 319774 292102
rect 319842 292046 319898 292102
rect 319718 291922 319774 291978
rect 319842 291922 319898 291978
rect 350438 292294 350494 292350
rect 350562 292294 350618 292350
rect 350438 292170 350494 292226
rect 350562 292170 350618 292226
rect 350438 292046 350494 292102
rect 350562 292046 350618 292102
rect 350438 291922 350494 291978
rect 350562 291922 350618 291978
rect 381158 292294 381214 292350
rect 381282 292294 381338 292350
rect 381158 292170 381214 292226
rect 381282 292170 381338 292226
rect 381158 292046 381214 292102
rect 381282 292046 381338 292102
rect 381158 291922 381214 291978
rect 381282 291922 381338 291978
rect 411878 292294 411934 292350
rect 412002 292294 412058 292350
rect 411878 292170 411934 292226
rect 412002 292170 412058 292226
rect 411878 292046 411934 292102
rect 412002 292046 412058 292102
rect 411878 291922 411934 291978
rect 412002 291922 412058 291978
rect 442598 292294 442654 292350
rect 442722 292294 442778 292350
rect 442598 292170 442654 292226
rect 442722 292170 442778 292226
rect 442598 292046 442654 292102
rect 442722 292046 442778 292102
rect 442598 291922 442654 291978
rect 442722 291922 442778 291978
rect 473318 292294 473374 292350
rect 473442 292294 473498 292350
rect 473318 292170 473374 292226
rect 473442 292170 473498 292226
rect 473318 292046 473374 292102
rect 473442 292046 473498 292102
rect 473318 291922 473374 291978
rect 473442 291922 473498 291978
rect 504038 292294 504094 292350
rect 504162 292294 504218 292350
rect 504038 292170 504094 292226
rect 504162 292170 504218 292226
rect 504038 292046 504094 292102
rect 504162 292046 504218 292102
rect 504038 291922 504094 291978
rect 504162 291922 504218 291978
rect 534758 292294 534814 292350
rect 534882 292294 534938 292350
rect 534758 292170 534814 292226
rect 534882 292170 534938 292226
rect 534758 292046 534814 292102
rect 534882 292046 534938 292102
rect 534758 291922 534814 291978
rect 534882 291922 534938 291978
rect 565478 292294 565534 292350
rect 565602 292294 565658 292350
rect 565478 292170 565534 292226
rect 565602 292170 565658 292226
rect 565478 292046 565534 292102
rect 565602 292046 565658 292102
rect 565478 291922 565534 291978
rect 565602 291922 565658 291978
rect 27878 280294 27934 280350
rect 28002 280294 28058 280350
rect 27878 280170 27934 280226
rect 28002 280170 28058 280226
rect 27878 280046 27934 280102
rect 28002 280046 28058 280102
rect 27878 279922 27934 279978
rect 28002 279922 28058 279978
rect 58598 280294 58654 280350
rect 58722 280294 58778 280350
rect 58598 280170 58654 280226
rect 58722 280170 58778 280226
rect 58598 280046 58654 280102
rect 58722 280046 58778 280102
rect 58598 279922 58654 279978
rect 58722 279922 58778 279978
rect 89318 280294 89374 280350
rect 89442 280294 89498 280350
rect 89318 280170 89374 280226
rect 89442 280170 89498 280226
rect 89318 280046 89374 280102
rect 89442 280046 89498 280102
rect 89318 279922 89374 279978
rect 89442 279922 89498 279978
rect 120038 280294 120094 280350
rect 120162 280294 120218 280350
rect 120038 280170 120094 280226
rect 120162 280170 120218 280226
rect 120038 280046 120094 280102
rect 120162 280046 120218 280102
rect 120038 279922 120094 279978
rect 120162 279922 120218 279978
rect 150758 280294 150814 280350
rect 150882 280294 150938 280350
rect 150758 280170 150814 280226
rect 150882 280170 150938 280226
rect 150758 280046 150814 280102
rect 150882 280046 150938 280102
rect 150758 279922 150814 279978
rect 150882 279922 150938 279978
rect 181478 280294 181534 280350
rect 181602 280294 181658 280350
rect 181478 280170 181534 280226
rect 181602 280170 181658 280226
rect 181478 280046 181534 280102
rect 181602 280046 181658 280102
rect 181478 279922 181534 279978
rect 181602 279922 181658 279978
rect 212198 280294 212254 280350
rect 212322 280294 212378 280350
rect 212198 280170 212254 280226
rect 212322 280170 212378 280226
rect 212198 280046 212254 280102
rect 212322 280046 212378 280102
rect 212198 279922 212254 279978
rect 212322 279922 212378 279978
rect 242918 280294 242974 280350
rect 243042 280294 243098 280350
rect 242918 280170 242974 280226
rect 243042 280170 243098 280226
rect 242918 280046 242974 280102
rect 243042 280046 243098 280102
rect 242918 279922 242974 279978
rect 243042 279922 243098 279978
rect 273638 280294 273694 280350
rect 273762 280294 273818 280350
rect 273638 280170 273694 280226
rect 273762 280170 273818 280226
rect 273638 280046 273694 280102
rect 273762 280046 273818 280102
rect 273638 279922 273694 279978
rect 273762 279922 273818 279978
rect 304358 280294 304414 280350
rect 304482 280294 304538 280350
rect 304358 280170 304414 280226
rect 304482 280170 304538 280226
rect 304358 280046 304414 280102
rect 304482 280046 304538 280102
rect 304358 279922 304414 279978
rect 304482 279922 304538 279978
rect 335078 280294 335134 280350
rect 335202 280294 335258 280350
rect 335078 280170 335134 280226
rect 335202 280170 335258 280226
rect 335078 280046 335134 280102
rect 335202 280046 335258 280102
rect 335078 279922 335134 279978
rect 335202 279922 335258 279978
rect 365798 280294 365854 280350
rect 365922 280294 365978 280350
rect 365798 280170 365854 280226
rect 365922 280170 365978 280226
rect 365798 280046 365854 280102
rect 365922 280046 365978 280102
rect 365798 279922 365854 279978
rect 365922 279922 365978 279978
rect 396518 280294 396574 280350
rect 396642 280294 396698 280350
rect 396518 280170 396574 280226
rect 396642 280170 396698 280226
rect 396518 280046 396574 280102
rect 396642 280046 396698 280102
rect 396518 279922 396574 279978
rect 396642 279922 396698 279978
rect 427238 280294 427294 280350
rect 427362 280294 427418 280350
rect 427238 280170 427294 280226
rect 427362 280170 427418 280226
rect 427238 280046 427294 280102
rect 427362 280046 427418 280102
rect 427238 279922 427294 279978
rect 427362 279922 427418 279978
rect 457958 280294 458014 280350
rect 458082 280294 458138 280350
rect 457958 280170 458014 280226
rect 458082 280170 458138 280226
rect 457958 280046 458014 280102
rect 458082 280046 458138 280102
rect 457958 279922 458014 279978
rect 458082 279922 458138 279978
rect 488678 280294 488734 280350
rect 488802 280294 488858 280350
rect 488678 280170 488734 280226
rect 488802 280170 488858 280226
rect 488678 280046 488734 280102
rect 488802 280046 488858 280102
rect 488678 279922 488734 279978
rect 488802 279922 488858 279978
rect 519398 280294 519454 280350
rect 519522 280294 519578 280350
rect 519398 280170 519454 280226
rect 519522 280170 519578 280226
rect 519398 280046 519454 280102
rect 519522 280046 519578 280102
rect 519398 279922 519454 279978
rect 519522 279922 519578 279978
rect 550118 280294 550174 280350
rect 550242 280294 550298 280350
rect 550118 280170 550174 280226
rect 550242 280170 550298 280226
rect 550118 280046 550174 280102
rect 550242 280046 550298 280102
rect 550118 279922 550174 279978
rect 550242 279922 550298 279978
rect 592914 352294 592970 352350
rect 593038 352294 593094 352350
rect 593162 352294 593218 352350
rect 593286 352294 593342 352350
rect 592914 352170 592970 352226
rect 593038 352170 593094 352226
rect 593162 352170 593218 352226
rect 593286 352170 593342 352226
rect 592914 352046 592970 352102
rect 593038 352046 593094 352102
rect 593162 352046 593218 352102
rect 593286 352046 593342 352102
rect 592914 351922 592970 351978
rect 593038 351922 593094 351978
rect 593162 351922 593218 351978
rect 593286 351922 593342 351978
rect 589194 328294 589250 328350
rect 589318 328294 589374 328350
rect 589442 328294 589498 328350
rect 589566 328294 589622 328350
rect 589194 328170 589250 328226
rect 589318 328170 589374 328226
rect 589442 328170 589498 328226
rect 589566 328170 589622 328226
rect 589194 328046 589250 328102
rect 589318 328046 589374 328102
rect 589442 328046 589498 328102
rect 589566 328046 589622 328102
rect 589194 327922 589250 327978
rect 589318 327922 589374 327978
rect 589442 327922 589498 327978
rect 589566 327922 589622 327978
rect 589194 310294 589250 310350
rect 589318 310294 589374 310350
rect 589442 310294 589498 310350
rect 589566 310294 589622 310350
rect 589194 310170 589250 310226
rect 589318 310170 589374 310226
rect 589442 310170 589498 310226
rect 589566 310170 589622 310226
rect 589194 310046 589250 310102
rect 589318 310046 589374 310102
rect 589442 310046 589498 310102
rect 589566 310046 589622 310102
rect 589194 309922 589250 309978
rect 589318 309922 589374 309978
rect 589442 309922 589498 309978
rect 589566 309922 589622 309978
rect 592914 334294 592970 334350
rect 593038 334294 593094 334350
rect 593162 334294 593218 334350
rect 593286 334294 593342 334350
rect 592914 334170 592970 334226
rect 593038 334170 593094 334226
rect 593162 334170 593218 334226
rect 593286 334170 593342 334226
rect 592914 334046 592970 334102
rect 593038 334046 593094 334102
rect 593162 334046 593218 334102
rect 593286 334046 593342 334102
rect 592914 333922 592970 333978
rect 593038 333922 593094 333978
rect 593162 333922 593218 333978
rect 593286 333922 593342 333978
rect 592914 316294 592970 316350
rect 593038 316294 593094 316350
rect 593162 316294 593218 316350
rect 593286 316294 593342 316350
rect 592914 316170 592970 316226
rect 593038 316170 593094 316226
rect 593162 316170 593218 316226
rect 593286 316170 593342 316226
rect 592914 316046 592970 316102
rect 593038 316046 593094 316102
rect 593162 316046 593218 316102
rect 593286 316046 593342 316102
rect 592914 315922 592970 315978
rect 593038 315922 593094 315978
rect 593162 315922 593218 315978
rect 593286 315922 593342 315978
rect 592914 298294 592970 298350
rect 593038 298294 593094 298350
rect 593162 298294 593218 298350
rect 593286 298294 593342 298350
rect 592914 298170 592970 298226
rect 593038 298170 593094 298226
rect 593162 298170 593218 298226
rect 593286 298170 593342 298226
rect 592914 298046 592970 298102
rect 593038 298046 593094 298102
rect 593162 298046 593218 298102
rect 593286 298046 593342 298102
rect 592914 297922 592970 297978
rect 593038 297922 593094 297978
rect 593162 297922 593218 297978
rect 593286 297922 593342 297978
rect 589194 292294 589250 292350
rect 589318 292294 589374 292350
rect 589442 292294 589498 292350
rect 589566 292294 589622 292350
rect 589194 292170 589250 292226
rect 589318 292170 589374 292226
rect 589442 292170 589498 292226
rect 589566 292170 589622 292226
rect 589194 292046 589250 292102
rect 589318 292046 589374 292102
rect 589442 292046 589498 292102
rect 589566 292046 589622 292102
rect 589194 291922 589250 291978
rect 589318 291922 589374 291978
rect 589442 291922 589498 291978
rect 589566 291922 589622 291978
rect 5514 274294 5570 274350
rect 5638 274294 5694 274350
rect 5762 274294 5818 274350
rect 5886 274294 5942 274350
rect 5514 274170 5570 274226
rect 5638 274170 5694 274226
rect 5762 274170 5818 274226
rect 5886 274170 5942 274226
rect 5514 274046 5570 274102
rect 5638 274046 5694 274102
rect 5762 274046 5818 274102
rect 5886 274046 5942 274102
rect 5514 273922 5570 273978
rect 5638 273922 5694 273978
rect 5762 273922 5818 273978
rect 5886 273922 5942 273978
rect -860 256294 -804 256350
rect -736 256294 -680 256350
rect -612 256294 -556 256350
rect -488 256294 -432 256350
rect -860 256170 -804 256226
rect -736 256170 -680 256226
rect -612 256170 -556 256226
rect -488 256170 -432 256226
rect -860 256046 -804 256102
rect -736 256046 -680 256102
rect -612 256046 -556 256102
rect -488 256046 -432 256102
rect -860 255922 -804 255978
rect -736 255922 -680 255978
rect -612 255922 -556 255978
rect -488 255922 -432 255978
rect -860 238294 -804 238350
rect -736 238294 -680 238350
rect -612 238294 -556 238350
rect -488 238294 -432 238350
rect -860 238170 -804 238226
rect -736 238170 -680 238226
rect -612 238170 -556 238226
rect -488 238170 -432 238226
rect -860 238046 -804 238102
rect -736 238046 -680 238102
rect -612 238046 -556 238102
rect -488 238046 -432 238102
rect -860 237922 -804 237978
rect -736 237922 -680 237978
rect -612 237922 -556 237978
rect -488 237922 -432 237978
rect 12518 274294 12574 274350
rect 12642 274294 12698 274350
rect 12518 274170 12574 274226
rect 12642 274170 12698 274226
rect 12518 274046 12574 274102
rect 12642 274046 12698 274102
rect 12518 273922 12574 273978
rect 12642 273922 12698 273978
rect 43238 274294 43294 274350
rect 43362 274294 43418 274350
rect 43238 274170 43294 274226
rect 43362 274170 43418 274226
rect 43238 274046 43294 274102
rect 43362 274046 43418 274102
rect 43238 273922 43294 273978
rect 43362 273922 43418 273978
rect 73958 274294 74014 274350
rect 74082 274294 74138 274350
rect 73958 274170 74014 274226
rect 74082 274170 74138 274226
rect 73958 274046 74014 274102
rect 74082 274046 74138 274102
rect 73958 273922 74014 273978
rect 74082 273922 74138 273978
rect 104678 274294 104734 274350
rect 104802 274294 104858 274350
rect 104678 274170 104734 274226
rect 104802 274170 104858 274226
rect 104678 274046 104734 274102
rect 104802 274046 104858 274102
rect 104678 273922 104734 273978
rect 104802 273922 104858 273978
rect 135398 274294 135454 274350
rect 135522 274294 135578 274350
rect 135398 274170 135454 274226
rect 135522 274170 135578 274226
rect 135398 274046 135454 274102
rect 135522 274046 135578 274102
rect 135398 273922 135454 273978
rect 135522 273922 135578 273978
rect 166118 274294 166174 274350
rect 166242 274294 166298 274350
rect 166118 274170 166174 274226
rect 166242 274170 166298 274226
rect 166118 274046 166174 274102
rect 166242 274046 166298 274102
rect 166118 273922 166174 273978
rect 166242 273922 166298 273978
rect 196838 274294 196894 274350
rect 196962 274294 197018 274350
rect 196838 274170 196894 274226
rect 196962 274170 197018 274226
rect 196838 274046 196894 274102
rect 196962 274046 197018 274102
rect 196838 273922 196894 273978
rect 196962 273922 197018 273978
rect 227558 274294 227614 274350
rect 227682 274294 227738 274350
rect 227558 274170 227614 274226
rect 227682 274170 227738 274226
rect 227558 274046 227614 274102
rect 227682 274046 227738 274102
rect 227558 273922 227614 273978
rect 227682 273922 227738 273978
rect 258278 274294 258334 274350
rect 258402 274294 258458 274350
rect 258278 274170 258334 274226
rect 258402 274170 258458 274226
rect 258278 274046 258334 274102
rect 258402 274046 258458 274102
rect 258278 273922 258334 273978
rect 258402 273922 258458 273978
rect 288998 274294 289054 274350
rect 289122 274294 289178 274350
rect 288998 274170 289054 274226
rect 289122 274170 289178 274226
rect 288998 274046 289054 274102
rect 289122 274046 289178 274102
rect 288998 273922 289054 273978
rect 289122 273922 289178 273978
rect 319718 274294 319774 274350
rect 319842 274294 319898 274350
rect 319718 274170 319774 274226
rect 319842 274170 319898 274226
rect 319718 274046 319774 274102
rect 319842 274046 319898 274102
rect 319718 273922 319774 273978
rect 319842 273922 319898 273978
rect 350438 274294 350494 274350
rect 350562 274294 350618 274350
rect 350438 274170 350494 274226
rect 350562 274170 350618 274226
rect 350438 274046 350494 274102
rect 350562 274046 350618 274102
rect 350438 273922 350494 273978
rect 350562 273922 350618 273978
rect 381158 274294 381214 274350
rect 381282 274294 381338 274350
rect 381158 274170 381214 274226
rect 381282 274170 381338 274226
rect 381158 274046 381214 274102
rect 381282 274046 381338 274102
rect 381158 273922 381214 273978
rect 381282 273922 381338 273978
rect 411878 274294 411934 274350
rect 412002 274294 412058 274350
rect 411878 274170 411934 274226
rect 412002 274170 412058 274226
rect 411878 274046 411934 274102
rect 412002 274046 412058 274102
rect 411878 273922 411934 273978
rect 412002 273922 412058 273978
rect 442598 274294 442654 274350
rect 442722 274294 442778 274350
rect 442598 274170 442654 274226
rect 442722 274170 442778 274226
rect 442598 274046 442654 274102
rect 442722 274046 442778 274102
rect 442598 273922 442654 273978
rect 442722 273922 442778 273978
rect 473318 274294 473374 274350
rect 473442 274294 473498 274350
rect 473318 274170 473374 274226
rect 473442 274170 473498 274226
rect 473318 274046 473374 274102
rect 473442 274046 473498 274102
rect 473318 273922 473374 273978
rect 473442 273922 473498 273978
rect 504038 274294 504094 274350
rect 504162 274294 504218 274350
rect 504038 274170 504094 274226
rect 504162 274170 504218 274226
rect 504038 274046 504094 274102
rect 504162 274046 504218 274102
rect 504038 273922 504094 273978
rect 504162 273922 504218 273978
rect 534758 274294 534814 274350
rect 534882 274294 534938 274350
rect 534758 274170 534814 274226
rect 534882 274170 534938 274226
rect 534758 274046 534814 274102
rect 534882 274046 534938 274102
rect 534758 273922 534814 273978
rect 534882 273922 534938 273978
rect 565478 274294 565534 274350
rect 565602 274294 565658 274350
rect 565478 274170 565534 274226
rect 565602 274170 565658 274226
rect 565478 274046 565534 274102
rect 565602 274046 565658 274102
rect 565478 273922 565534 273978
rect 565602 273922 565658 273978
rect 5514 256294 5570 256350
rect 5638 256294 5694 256350
rect 5762 256294 5818 256350
rect 5886 256294 5942 256350
rect 5514 256170 5570 256226
rect 5638 256170 5694 256226
rect 5762 256170 5818 256226
rect 5886 256170 5942 256226
rect 5514 256046 5570 256102
rect 5638 256046 5694 256102
rect 5762 256046 5818 256102
rect 5886 256046 5942 256102
rect 5514 255922 5570 255978
rect 5638 255922 5694 255978
rect 5762 255922 5818 255978
rect 5886 255922 5942 255978
rect 27878 262294 27934 262350
rect 28002 262294 28058 262350
rect 27878 262170 27934 262226
rect 28002 262170 28058 262226
rect 27878 262046 27934 262102
rect 28002 262046 28058 262102
rect 27878 261922 27934 261978
rect 28002 261922 28058 261978
rect 58598 262294 58654 262350
rect 58722 262294 58778 262350
rect 58598 262170 58654 262226
rect 58722 262170 58778 262226
rect 58598 262046 58654 262102
rect 58722 262046 58778 262102
rect 58598 261922 58654 261978
rect 58722 261922 58778 261978
rect 89318 262294 89374 262350
rect 89442 262294 89498 262350
rect 89318 262170 89374 262226
rect 89442 262170 89498 262226
rect 89318 262046 89374 262102
rect 89442 262046 89498 262102
rect 89318 261922 89374 261978
rect 89442 261922 89498 261978
rect 120038 262294 120094 262350
rect 120162 262294 120218 262350
rect 120038 262170 120094 262226
rect 120162 262170 120218 262226
rect 120038 262046 120094 262102
rect 120162 262046 120218 262102
rect 120038 261922 120094 261978
rect 120162 261922 120218 261978
rect 150758 262294 150814 262350
rect 150882 262294 150938 262350
rect 150758 262170 150814 262226
rect 150882 262170 150938 262226
rect 150758 262046 150814 262102
rect 150882 262046 150938 262102
rect 150758 261922 150814 261978
rect 150882 261922 150938 261978
rect 181478 262294 181534 262350
rect 181602 262294 181658 262350
rect 181478 262170 181534 262226
rect 181602 262170 181658 262226
rect 181478 262046 181534 262102
rect 181602 262046 181658 262102
rect 181478 261922 181534 261978
rect 181602 261922 181658 261978
rect 212198 262294 212254 262350
rect 212322 262294 212378 262350
rect 212198 262170 212254 262226
rect 212322 262170 212378 262226
rect 212198 262046 212254 262102
rect 212322 262046 212378 262102
rect 212198 261922 212254 261978
rect 212322 261922 212378 261978
rect 242918 262294 242974 262350
rect 243042 262294 243098 262350
rect 242918 262170 242974 262226
rect 243042 262170 243098 262226
rect 242918 262046 242974 262102
rect 243042 262046 243098 262102
rect 242918 261922 242974 261978
rect 243042 261922 243098 261978
rect 273638 262294 273694 262350
rect 273762 262294 273818 262350
rect 273638 262170 273694 262226
rect 273762 262170 273818 262226
rect 273638 262046 273694 262102
rect 273762 262046 273818 262102
rect 273638 261922 273694 261978
rect 273762 261922 273818 261978
rect 304358 262294 304414 262350
rect 304482 262294 304538 262350
rect 304358 262170 304414 262226
rect 304482 262170 304538 262226
rect 304358 262046 304414 262102
rect 304482 262046 304538 262102
rect 304358 261922 304414 261978
rect 304482 261922 304538 261978
rect 335078 262294 335134 262350
rect 335202 262294 335258 262350
rect 335078 262170 335134 262226
rect 335202 262170 335258 262226
rect 335078 262046 335134 262102
rect 335202 262046 335258 262102
rect 335078 261922 335134 261978
rect 335202 261922 335258 261978
rect 365798 262294 365854 262350
rect 365922 262294 365978 262350
rect 365798 262170 365854 262226
rect 365922 262170 365978 262226
rect 365798 262046 365854 262102
rect 365922 262046 365978 262102
rect 365798 261922 365854 261978
rect 365922 261922 365978 261978
rect 396518 262294 396574 262350
rect 396642 262294 396698 262350
rect 396518 262170 396574 262226
rect 396642 262170 396698 262226
rect 396518 262046 396574 262102
rect 396642 262046 396698 262102
rect 396518 261922 396574 261978
rect 396642 261922 396698 261978
rect 427238 262294 427294 262350
rect 427362 262294 427418 262350
rect 427238 262170 427294 262226
rect 427362 262170 427418 262226
rect 427238 262046 427294 262102
rect 427362 262046 427418 262102
rect 427238 261922 427294 261978
rect 427362 261922 427418 261978
rect 457958 262294 458014 262350
rect 458082 262294 458138 262350
rect 457958 262170 458014 262226
rect 458082 262170 458138 262226
rect 457958 262046 458014 262102
rect 458082 262046 458138 262102
rect 457958 261922 458014 261978
rect 458082 261922 458138 261978
rect 488678 262294 488734 262350
rect 488802 262294 488858 262350
rect 488678 262170 488734 262226
rect 488802 262170 488858 262226
rect 488678 262046 488734 262102
rect 488802 262046 488858 262102
rect 488678 261922 488734 261978
rect 488802 261922 488858 261978
rect 519398 262294 519454 262350
rect 519522 262294 519578 262350
rect 519398 262170 519454 262226
rect 519522 262170 519578 262226
rect 519398 262046 519454 262102
rect 519522 262046 519578 262102
rect 519398 261922 519454 261978
rect 519522 261922 519578 261978
rect 550118 262294 550174 262350
rect 550242 262294 550298 262350
rect 550118 262170 550174 262226
rect 550242 262170 550298 262226
rect 550118 262046 550174 262102
rect 550242 262046 550298 262102
rect 550118 261922 550174 261978
rect 550242 261922 550298 261978
rect 12518 256294 12574 256350
rect 12642 256294 12698 256350
rect 12518 256170 12574 256226
rect 12642 256170 12698 256226
rect 12518 256046 12574 256102
rect 12642 256046 12698 256102
rect 12518 255922 12574 255978
rect 12642 255922 12698 255978
rect 43238 256294 43294 256350
rect 43362 256294 43418 256350
rect 43238 256170 43294 256226
rect 43362 256170 43418 256226
rect 43238 256046 43294 256102
rect 43362 256046 43418 256102
rect 43238 255922 43294 255978
rect 43362 255922 43418 255978
rect 73958 256294 74014 256350
rect 74082 256294 74138 256350
rect 73958 256170 74014 256226
rect 74082 256170 74138 256226
rect 73958 256046 74014 256102
rect 74082 256046 74138 256102
rect 73958 255922 74014 255978
rect 74082 255922 74138 255978
rect 104678 256294 104734 256350
rect 104802 256294 104858 256350
rect 104678 256170 104734 256226
rect 104802 256170 104858 256226
rect 104678 256046 104734 256102
rect 104802 256046 104858 256102
rect 104678 255922 104734 255978
rect 104802 255922 104858 255978
rect 135398 256294 135454 256350
rect 135522 256294 135578 256350
rect 135398 256170 135454 256226
rect 135522 256170 135578 256226
rect 135398 256046 135454 256102
rect 135522 256046 135578 256102
rect 135398 255922 135454 255978
rect 135522 255922 135578 255978
rect 166118 256294 166174 256350
rect 166242 256294 166298 256350
rect 166118 256170 166174 256226
rect 166242 256170 166298 256226
rect 166118 256046 166174 256102
rect 166242 256046 166298 256102
rect 166118 255922 166174 255978
rect 166242 255922 166298 255978
rect 196838 256294 196894 256350
rect 196962 256294 197018 256350
rect 196838 256170 196894 256226
rect 196962 256170 197018 256226
rect 196838 256046 196894 256102
rect 196962 256046 197018 256102
rect 196838 255922 196894 255978
rect 196962 255922 197018 255978
rect 227558 256294 227614 256350
rect 227682 256294 227738 256350
rect 227558 256170 227614 256226
rect 227682 256170 227738 256226
rect 227558 256046 227614 256102
rect 227682 256046 227738 256102
rect 227558 255922 227614 255978
rect 227682 255922 227738 255978
rect 258278 256294 258334 256350
rect 258402 256294 258458 256350
rect 258278 256170 258334 256226
rect 258402 256170 258458 256226
rect 258278 256046 258334 256102
rect 258402 256046 258458 256102
rect 258278 255922 258334 255978
rect 258402 255922 258458 255978
rect 288998 256294 289054 256350
rect 289122 256294 289178 256350
rect 288998 256170 289054 256226
rect 289122 256170 289178 256226
rect 288998 256046 289054 256102
rect 289122 256046 289178 256102
rect 288998 255922 289054 255978
rect 289122 255922 289178 255978
rect 319718 256294 319774 256350
rect 319842 256294 319898 256350
rect 319718 256170 319774 256226
rect 319842 256170 319898 256226
rect 319718 256046 319774 256102
rect 319842 256046 319898 256102
rect 319718 255922 319774 255978
rect 319842 255922 319898 255978
rect 350438 256294 350494 256350
rect 350562 256294 350618 256350
rect 350438 256170 350494 256226
rect 350562 256170 350618 256226
rect 350438 256046 350494 256102
rect 350562 256046 350618 256102
rect 350438 255922 350494 255978
rect 350562 255922 350618 255978
rect 381158 256294 381214 256350
rect 381282 256294 381338 256350
rect 381158 256170 381214 256226
rect 381282 256170 381338 256226
rect 381158 256046 381214 256102
rect 381282 256046 381338 256102
rect 381158 255922 381214 255978
rect 381282 255922 381338 255978
rect 411878 256294 411934 256350
rect 412002 256294 412058 256350
rect 411878 256170 411934 256226
rect 412002 256170 412058 256226
rect 411878 256046 411934 256102
rect 412002 256046 412058 256102
rect 411878 255922 411934 255978
rect 412002 255922 412058 255978
rect 442598 256294 442654 256350
rect 442722 256294 442778 256350
rect 442598 256170 442654 256226
rect 442722 256170 442778 256226
rect 442598 256046 442654 256102
rect 442722 256046 442778 256102
rect 442598 255922 442654 255978
rect 442722 255922 442778 255978
rect 473318 256294 473374 256350
rect 473442 256294 473498 256350
rect 473318 256170 473374 256226
rect 473442 256170 473498 256226
rect 473318 256046 473374 256102
rect 473442 256046 473498 256102
rect 473318 255922 473374 255978
rect 473442 255922 473498 255978
rect 504038 256294 504094 256350
rect 504162 256294 504218 256350
rect 504038 256170 504094 256226
rect 504162 256170 504218 256226
rect 504038 256046 504094 256102
rect 504162 256046 504218 256102
rect 504038 255922 504094 255978
rect 504162 255922 504218 255978
rect 534758 256294 534814 256350
rect 534882 256294 534938 256350
rect 534758 256170 534814 256226
rect 534882 256170 534938 256226
rect 534758 256046 534814 256102
rect 534882 256046 534938 256102
rect 534758 255922 534814 255978
rect 534882 255922 534938 255978
rect 565478 256294 565534 256350
rect 565602 256294 565658 256350
rect 565478 256170 565534 256226
rect 565602 256170 565658 256226
rect 565478 256046 565534 256102
rect 565602 256046 565658 256102
rect 565478 255922 565534 255978
rect 565602 255922 565658 255978
rect 5514 238294 5570 238350
rect 5638 238294 5694 238350
rect 5762 238294 5818 238350
rect 5886 238294 5942 238350
rect 5514 238170 5570 238226
rect 5638 238170 5694 238226
rect 5762 238170 5818 238226
rect 5886 238170 5942 238226
rect 5514 238046 5570 238102
rect 5638 238046 5694 238102
rect 5762 238046 5818 238102
rect 5886 238046 5942 238102
rect 5514 237922 5570 237978
rect 5638 237922 5694 237978
rect 5762 237922 5818 237978
rect 5886 237922 5942 237978
rect -860 220294 -804 220350
rect -736 220294 -680 220350
rect -612 220294 -556 220350
rect -488 220294 -432 220350
rect -860 220170 -804 220226
rect -736 220170 -680 220226
rect -612 220170 -556 220226
rect -488 220170 -432 220226
rect -860 220046 -804 220102
rect -736 220046 -680 220102
rect -612 220046 -556 220102
rect -488 220046 -432 220102
rect -860 219922 -804 219978
rect -736 219922 -680 219978
rect -612 219922 -556 219978
rect -488 219922 -432 219978
rect 27878 244294 27934 244350
rect 28002 244294 28058 244350
rect 27878 244170 27934 244226
rect 28002 244170 28058 244226
rect 27878 244046 27934 244102
rect 28002 244046 28058 244102
rect 27878 243922 27934 243978
rect 28002 243922 28058 243978
rect 58598 244294 58654 244350
rect 58722 244294 58778 244350
rect 58598 244170 58654 244226
rect 58722 244170 58778 244226
rect 58598 244046 58654 244102
rect 58722 244046 58778 244102
rect 58598 243922 58654 243978
rect 58722 243922 58778 243978
rect 89318 244294 89374 244350
rect 89442 244294 89498 244350
rect 89318 244170 89374 244226
rect 89442 244170 89498 244226
rect 89318 244046 89374 244102
rect 89442 244046 89498 244102
rect 89318 243922 89374 243978
rect 89442 243922 89498 243978
rect 120038 244294 120094 244350
rect 120162 244294 120218 244350
rect 120038 244170 120094 244226
rect 120162 244170 120218 244226
rect 120038 244046 120094 244102
rect 120162 244046 120218 244102
rect 120038 243922 120094 243978
rect 120162 243922 120218 243978
rect 150758 244294 150814 244350
rect 150882 244294 150938 244350
rect 150758 244170 150814 244226
rect 150882 244170 150938 244226
rect 150758 244046 150814 244102
rect 150882 244046 150938 244102
rect 150758 243922 150814 243978
rect 150882 243922 150938 243978
rect 181478 244294 181534 244350
rect 181602 244294 181658 244350
rect 181478 244170 181534 244226
rect 181602 244170 181658 244226
rect 181478 244046 181534 244102
rect 181602 244046 181658 244102
rect 181478 243922 181534 243978
rect 181602 243922 181658 243978
rect 212198 244294 212254 244350
rect 212322 244294 212378 244350
rect 212198 244170 212254 244226
rect 212322 244170 212378 244226
rect 212198 244046 212254 244102
rect 212322 244046 212378 244102
rect 212198 243922 212254 243978
rect 212322 243922 212378 243978
rect 242918 244294 242974 244350
rect 243042 244294 243098 244350
rect 242918 244170 242974 244226
rect 243042 244170 243098 244226
rect 242918 244046 242974 244102
rect 243042 244046 243098 244102
rect 242918 243922 242974 243978
rect 243042 243922 243098 243978
rect 273638 244294 273694 244350
rect 273762 244294 273818 244350
rect 273638 244170 273694 244226
rect 273762 244170 273818 244226
rect 273638 244046 273694 244102
rect 273762 244046 273818 244102
rect 273638 243922 273694 243978
rect 273762 243922 273818 243978
rect 304358 244294 304414 244350
rect 304482 244294 304538 244350
rect 304358 244170 304414 244226
rect 304482 244170 304538 244226
rect 304358 244046 304414 244102
rect 304482 244046 304538 244102
rect 304358 243922 304414 243978
rect 304482 243922 304538 243978
rect 335078 244294 335134 244350
rect 335202 244294 335258 244350
rect 335078 244170 335134 244226
rect 335202 244170 335258 244226
rect 335078 244046 335134 244102
rect 335202 244046 335258 244102
rect 335078 243922 335134 243978
rect 335202 243922 335258 243978
rect 365798 244294 365854 244350
rect 365922 244294 365978 244350
rect 365798 244170 365854 244226
rect 365922 244170 365978 244226
rect 365798 244046 365854 244102
rect 365922 244046 365978 244102
rect 365798 243922 365854 243978
rect 365922 243922 365978 243978
rect 396518 244294 396574 244350
rect 396642 244294 396698 244350
rect 396518 244170 396574 244226
rect 396642 244170 396698 244226
rect 396518 244046 396574 244102
rect 396642 244046 396698 244102
rect 396518 243922 396574 243978
rect 396642 243922 396698 243978
rect 427238 244294 427294 244350
rect 427362 244294 427418 244350
rect 427238 244170 427294 244226
rect 427362 244170 427418 244226
rect 427238 244046 427294 244102
rect 427362 244046 427418 244102
rect 427238 243922 427294 243978
rect 427362 243922 427418 243978
rect 457958 244294 458014 244350
rect 458082 244294 458138 244350
rect 457958 244170 458014 244226
rect 458082 244170 458138 244226
rect 457958 244046 458014 244102
rect 458082 244046 458138 244102
rect 457958 243922 458014 243978
rect 458082 243922 458138 243978
rect 488678 244294 488734 244350
rect 488802 244294 488858 244350
rect 488678 244170 488734 244226
rect 488802 244170 488858 244226
rect 488678 244046 488734 244102
rect 488802 244046 488858 244102
rect 488678 243922 488734 243978
rect 488802 243922 488858 243978
rect 519398 244294 519454 244350
rect 519522 244294 519578 244350
rect 519398 244170 519454 244226
rect 519522 244170 519578 244226
rect 519398 244046 519454 244102
rect 519522 244046 519578 244102
rect 519398 243922 519454 243978
rect 519522 243922 519578 243978
rect 550118 244294 550174 244350
rect 550242 244294 550298 244350
rect 550118 244170 550174 244226
rect 550242 244170 550298 244226
rect 550118 244046 550174 244102
rect 550242 244046 550298 244102
rect 550118 243922 550174 243978
rect 550242 243922 550298 243978
rect 12518 238294 12574 238350
rect 12642 238294 12698 238350
rect 12518 238170 12574 238226
rect 12642 238170 12698 238226
rect 12518 238046 12574 238102
rect 12642 238046 12698 238102
rect 12518 237922 12574 237978
rect 12642 237922 12698 237978
rect 43238 238294 43294 238350
rect 43362 238294 43418 238350
rect 43238 238170 43294 238226
rect 43362 238170 43418 238226
rect 43238 238046 43294 238102
rect 43362 238046 43418 238102
rect 43238 237922 43294 237978
rect 43362 237922 43418 237978
rect 73958 238294 74014 238350
rect 74082 238294 74138 238350
rect 73958 238170 74014 238226
rect 74082 238170 74138 238226
rect 73958 238046 74014 238102
rect 74082 238046 74138 238102
rect 73958 237922 74014 237978
rect 74082 237922 74138 237978
rect 104678 238294 104734 238350
rect 104802 238294 104858 238350
rect 104678 238170 104734 238226
rect 104802 238170 104858 238226
rect 104678 238046 104734 238102
rect 104802 238046 104858 238102
rect 104678 237922 104734 237978
rect 104802 237922 104858 237978
rect 135398 238294 135454 238350
rect 135522 238294 135578 238350
rect 135398 238170 135454 238226
rect 135522 238170 135578 238226
rect 135398 238046 135454 238102
rect 135522 238046 135578 238102
rect 135398 237922 135454 237978
rect 135522 237922 135578 237978
rect 166118 238294 166174 238350
rect 166242 238294 166298 238350
rect 166118 238170 166174 238226
rect 166242 238170 166298 238226
rect 166118 238046 166174 238102
rect 166242 238046 166298 238102
rect 166118 237922 166174 237978
rect 166242 237922 166298 237978
rect 196838 238294 196894 238350
rect 196962 238294 197018 238350
rect 196838 238170 196894 238226
rect 196962 238170 197018 238226
rect 196838 238046 196894 238102
rect 196962 238046 197018 238102
rect 196838 237922 196894 237978
rect 196962 237922 197018 237978
rect 227558 238294 227614 238350
rect 227682 238294 227738 238350
rect 227558 238170 227614 238226
rect 227682 238170 227738 238226
rect 227558 238046 227614 238102
rect 227682 238046 227738 238102
rect 227558 237922 227614 237978
rect 227682 237922 227738 237978
rect 258278 238294 258334 238350
rect 258402 238294 258458 238350
rect 258278 238170 258334 238226
rect 258402 238170 258458 238226
rect 258278 238046 258334 238102
rect 258402 238046 258458 238102
rect 258278 237922 258334 237978
rect 258402 237922 258458 237978
rect 288998 238294 289054 238350
rect 289122 238294 289178 238350
rect 288998 238170 289054 238226
rect 289122 238170 289178 238226
rect 288998 238046 289054 238102
rect 289122 238046 289178 238102
rect 288998 237922 289054 237978
rect 289122 237922 289178 237978
rect 319718 238294 319774 238350
rect 319842 238294 319898 238350
rect 319718 238170 319774 238226
rect 319842 238170 319898 238226
rect 319718 238046 319774 238102
rect 319842 238046 319898 238102
rect 319718 237922 319774 237978
rect 319842 237922 319898 237978
rect 350438 238294 350494 238350
rect 350562 238294 350618 238350
rect 350438 238170 350494 238226
rect 350562 238170 350618 238226
rect 350438 238046 350494 238102
rect 350562 238046 350618 238102
rect 350438 237922 350494 237978
rect 350562 237922 350618 237978
rect 381158 238294 381214 238350
rect 381282 238294 381338 238350
rect 381158 238170 381214 238226
rect 381282 238170 381338 238226
rect 381158 238046 381214 238102
rect 381282 238046 381338 238102
rect 381158 237922 381214 237978
rect 381282 237922 381338 237978
rect 411878 238294 411934 238350
rect 412002 238294 412058 238350
rect 411878 238170 411934 238226
rect 412002 238170 412058 238226
rect 411878 238046 411934 238102
rect 412002 238046 412058 238102
rect 411878 237922 411934 237978
rect 412002 237922 412058 237978
rect 442598 238294 442654 238350
rect 442722 238294 442778 238350
rect 442598 238170 442654 238226
rect 442722 238170 442778 238226
rect 442598 238046 442654 238102
rect 442722 238046 442778 238102
rect 442598 237922 442654 237978
rect 442722 237922 442778 237978
rect 473318 238294 473374 238350
rect 473442 238294 473498 238350
rect 473318 238170 473374 238226
rect 473442 238170 473498 238226
rect 473318 238046 473374 238102
rect 473442 238046 473498 238102
rect 473318 237922 473374 237978
rect 473442 237922 473498 237978
rect 504038 238294 504094 238350
rect 504162 238294 504218 238350
rect 504038 238170 504094 238226
rect 504162 238170 504218 238226
rect 504038 238046 504094 238102
rect 504162 238046 504218 238102
rect 504038 237922 504094 237978
rect 504162 237922 504218 237978
rect 534758 238294 534814 238350
rect 534882 238294 534938 238350
rect 534758 238170 534814 238226
rect 534882 238170 534938 238226
rect 534758 238046 534814 238102
rect 534882 238046 534938 238102
rect 534758 237922 534814 237978
rect 534882 237922 534938 237978
rect 565478 238294 565534 238350
rect 565602 238294 565658 238350
rect 565478 238170 565534 238226
rect 565602 238170 565658 238226
rect 565478 238046 565534 238102
rect 565602 238046 565658 238102
rect 565478 237922 565534 237978
rect 565602 237922 565658 237978
rect 589194 274294 589250 274350
rect 589318 274294 589374 274350
rect 589442 274294 589498 274350
rect 589566 274294 589622 274350
rect 589194 274170 589250 274226
rect 589318 274170 589374 274226
rect 589442 274170 589498 274226
rect 589566 274170 589622 274226
rect 589194 274046 589250 274102
rect 589318 274046 589374 274102
rect 589442 274046 589498 274102
rect 589566 274046 589622 274102
rect 589194 273922 589250 273978
rect 589318 273922 589374 273978
rect 589442 273922 589498 273978
rect 589566 273922 589622 273978
rect 27878 226294 27934 226350
rect 28002 226294 28058 226350
rect 27878 226170 27934 226226
rect 28002 226170 28058 226226
rect 27878 226046 27934 226102
rect 28002 226046 28058 226102
rect 27878 225922 27934 225978
rect 28002 225922 28058 225978
rect 58598 226294 58654 226350
rect 58722 226294 58778 226350
rect 58598 226170 58654 226226
rect 58722 226170 58778 226226
rect 58598 226046 58654 226102
rect 58722 226046 58778 226102
rect 58598 225922 58654 225978
rect 58722 225922 58778 225978
rect 89318 226294 89374 226350
rect 89442 226294 89498 226350
rect 89318 226170 89374 226226
rect 89442 226170 89498 226226
rect 89318 226046 89374 226102
rect 89442 226046 89498 226102
rect 89318 225922 89374 225978
rect 89442 225922 89498 225978
rect 120038 226294 120094 226350
rect 120162 226294 120218 226350
rect 120038 226170 120094 226226
rect 120162 226170 120218 226226
rect 120038 226046 120094 226102
rect 120162 226046 120218 226102
rect 120038 225922 120094 225978
rect 120162 225922 120218 225978
rect 150758 226294 150814 226350
rect 150882 226294 150938 226350
rect 150758 226170 150814 226226
rect 150882 226170 150938 226226
rect 150758 226046 150814 226102
rect 150882 226046 150938 226102
rect 150758 225922 150814 225978
rect 150882 225922 150938 225978
rect 181478 226294 181534 226350
rect 181602 226294 181658 226350
rect 181478 226170 181534 226226
rect 181602 226170 181658 226226
rect 181478 226046 181534 226102
rect 181602 226046 181658 226102
rect 181478 225922 181534 225978
rect 181602 225922 181658 225978
rect 212198 226294 212254 226350
rect 212322 226294 212378 226350
rect 212198 226170 212254 226226
rect 212322 226170 212378 226226
rect 212198 226046 212254 226102
rect 212322 226046 212378 226102
rect 212198 225922 212254 225978
rect 212322 225922 212378 225978
rect 242918 226294 242974 226350
rect 243042 226294 243098 226350
rect 242918 226170 242974 226226
rect 243042 226170 243098 226226
rect 242918 226046 242974 226102
rect 243042 226046 243098 226102
rect 242918 225922 242974 225978
rect 243042 225922 243098 225978
rect 273638 226294 273694 226350
rect 273762 226294 273818 226350
rect 273638 226170 273694 226226
rect 273762 226170 273818 226226
rect 273638 226046 273694 226102
rect 273762 226046 273818 226102
rect 273638 225922 273694 225978
rect 273762 225922 273818 225978
rect 304358 226294 304414 226350
rect 304482 226294 304538 226350
rect 304358 226170 304414 226226
rect 304482 226170 304538 226226
rect 304358 226046 304414 226102
rect 304482 226046 304538 226102
rect 304358 225922 304414 225978
rect 304482 225922 304538 225978
rect 335078 226294 335134 226350
rect 335202 226294 335258 226350
rect 335078 226170 335134 226226
rect 335202 226170 335258 226226
rect 335078 226046 335134 226102
rect 335202 226046 335258 226102
rect 335078 225922 335134 225978
rect 335202 225922 335258 225978
rect 365798 226294 365854 226350
rect 365922 226294 365978 226350
rect 365798 226170 365854 226226
rect 365922 226170 365978 226226
rect 365798 226046 365854 226102
rect 365922 226046 365978 226102
rect 365798 225922 365854 225978
rect 365922 225922 365978 225978
rect 396518 226294 396574 226350
rect 396642 226294 396698 226350
rect 396518 226170 396574 226226
rect 396642 226170 396698 226226
rect 396518 226046 396574 226102
rect 396642 226046 396698 226102
rect 396518 225922 396574 225978
rect 396642 225922 396698 225978
rect 427238 226294 427294 226350
rect 427362 226294 427418 226350
rect 427238 226170 427294 226226
rect 427362 226170 427418 226226
rect 427238 226046 427294 226102
rect 427362 226046 427418 226102
rect 427238 225922 427294 225978
rect 427362 225922 427418 225978
rect 457958 226294 458014 226350
rect 458082 226294 458138 226350
rect 457958 226170 458014 226226
rect 458082 226170 458138 226226
rect 457958 226046 458014 226102
rect 458082 226046 458138 226102
rect 457958 225922 458014 225978
rect 458082 225922 458138 225978
rect 488678 226294 488734 226350
rect 488802 226294 488858 226350
rect 488678 226170 488734 226226
rect 488802 226170 488858 226226
rect 488678 226046 488734 226102
rect 488802 226046 488858 226102
rect 488678 225922 488734 225978
rect 488802 225922 488858 225978
rect 519398 226294 519454 226350
rect 519522 226294 519578 226350
rect 519398 226170 519454 226226
rect 519522 226170 519578 226226
rect 519398 226046 519454 226102
rect 519522 226046 519578 226102
rect 519398 225922 519454 225978
rect 519522 225922 519578 225978
rect 550118 226294 550174 226350
rect 550242 226294 550298 226350
rect 550118 226170 550174 226226
rect 550242 226170 550298 226226
rect 550118 226046 550174 226102
rect 550242 226046 550298 226102
rect 550118 225922 550174 225978
rect 550242 225922 550298 225978
rect 5514 220294 5570 220350
rect 5638 220294 5694 220350
rect 5762 220294 5818 220350
rect 5886 220294 5942 220350
rect 12518 220294 12574 220350
rect 12642 220294 12698 220350
rect 5514 220170 5570 220226
rect 5638 220170 5694 220226
rect 5762 220170 5818 220226
rect 5886 220170 5942 220226
rect 5514 220046 5570 220102
rect 5638 220046 5694 220102
rect 5762 220046 5818 220102
rect 5886 220046 5942 220102
rect 5514 219922 5570 219978
rect 5638 219922 5694 219978
rect 5762 219922 5818 219978
rect 5886 219922 5942 219978
rect -860 202294 -804 202350
rect -736 202294 -680 202350
rect -612 202294 -556 202350
rect -488 202294 -432 202350
rect -860 202170 -804 202226
rect -736 202170 -680 202226
rect -612 202170 -556 202226
rect -488 202170 -432 202226
rect -860 202046 -804 202102
rect -736 202046 -680 202102
rect -612 202046 -556 202102
rect -488 202046 -432 202102
rect -860 201922 -804 201978
rect -736 201922 -680 201978
rect -612 201922 -556 201978
rect -488 201922 -432 201978
rect 12518 220170 12574 220226
rect 12642 220170 12698 220226
rect 12518 220046 12574 220102
rect 12642 220046 12698 220102
rect 12518 219922 12574 219978
rect 12642 219922 12698 219978
rect 43238 220294 43294 220350
rect 43362 220294 43418 220350
rect 43238 220170 43294 220226
rect 43362 220170 43418 220226
rect 43238 220046 43294 220102
rect 43362 220046 43418 220102
rect 43238 219922 43294 219978
rect 43362 219922 43418 219978
rect 73958 220294 74014 220350
rect 74082 220294 74138 220350
rect 73958 220170 74014 220226
rect 74082 220170 74138 220226
rect 73958 220046 74014 220102
rect 74082 220046 74138 220102
rect 73958 219922 74014 219978
rect 74082 219922 74138 219978
rect 104678 220294 104734 220350
rect 104802 220294 104858 220350
rect 104678 220170 104734 220226
rect 104802 220170 104858 220226
rect 104678 220046 104734 220102
rect 104802 220046 104858 220102
rect 104678 219922 104734 219978
rect 104802 219922 104858 219978
rect 135398 220294 135454 220350
rect 135522 220294 135578 220350
rect 135398 220170 135454 220226
rect 135522 220170 135578 220226
rect 135398 220046 135454 220102
rect 135522 220046 135578 220102
rect 135398 219922 135454 219978
rect 135522 219922 135578 219978
rect 166118 220294 166174 220350
rect 166242 220294 166298 220350
rect 166118 220170 166174 220226
rect 166242 220170 166298 220226
rect 166118 220046 166174 220102
rect 166242 220046 166298 220102
rect 166118 219922 166174 219978
rect 166242 219922 166298 219978
rect 196838 220294 196894 220350
rect 196962 220294 197018 220350
rect 196838 220170 196894 220226
rect 196962 220170 197018 220226
rect 196838 220046 196894 220102
rect 196962 220046 197018 220102
rect 196838 219922 196894 219978
rect 196962 219922 197018 219978
rect 227558 220294 227614 220350
rect 227682 220294 227738 220350
rect 227558 220170 227614 220226
rect 227682 220170 227738 220226
rect 227558 220046 227614 220102
rect 227682 220046 227738 220102
rect 227558 219922 227614 219978
rect 227682 219922 227738 219978
rect 258278 220294 258334 220350
rect 258402 220294 258458 220350
rect 258278 220170 258334 220226
rect 258402 220170 258458 220226
rect 258278 220046 258334 220102
rect 258402 220046 258458 220102
rect 258278 219922 258334 219978
rect 258402 219922 258458 219978
rect 288998 220294 289054 220350
rect 289122 220294 289178 220350
rect 288998 220170 289054 220226
rect 289122 220170 289178 220226
rect 288998 220046 289054 220102
rect 289122 220046 289178 220102
rect 288998 219922 289054 219978
rect 289122 219922 289178 219978
rect 319718 220294 319774 220350
rect 319842 220294 319898 220350
rect 319718 220170 319774 220226
rect 319842 220170 319898 220226
rect 319718 220046 319774 220102
rect 319842 220046 319898 220102
rect 319718 219922 319774 219978
rect 319842 219922 319898 219978
rect 350438 220294 350494 220350
rect 350562 220294 350618 220350
rect 350438 220170 350494 220226
rect 350562 220170 350618 220226
rect 350438 220046 350494 220102
rect 350562 220046 350618 220102
rect 350438 219922 350494 219978
rect 350562 219922 350618 219978
rect 381158 220294 381214 220350
rect 381282 220294 381338 220350
rect 381158 220170 381214 220226
rect 381282 220170 381338 220226
rect 381158 220046 381214 220102
rect 381282 220046 381338 220102
rect 381158 219922 381214 219978
rect 381282 219922 381338 219978
rect 411878 220294 411934 220350
rect 412002 220294 412058 220350
rect 411878 220170 411934 220226
rect 412002 220170 412058 220226
rect 411878 220046 411934 220102
rect 412002 220046 412058 220102
rect 411878 219922 411934 219978
rect 412002 219922 412058 219978
rect 442598 220294 442654 220350
rect 442722 220294 442778 220350
rect 442598 220170 442654 220226
rect 442722 220170 442778 220226
rect 442598 220046 442654 220102
rect 442722 220046 442778 220102
rect 442598 219922 442654 219978
rect 442722 219922 442778 219978
rect 473318 220294 473374 220350
rect 473442 220294 473498 220350
rect 473318 220170 473374 220226
rect 473442 220170 473498 220226
rect 473318 220046 473374 220102
rect 473442 220046 473498 220102
rect 473318 219922 473374 219978
rect 473442 219922 473498 219978
rect 504038 220294 504094 220350
rect 504162 220294 504218 220350
rect 504038 220170 504094 220226
rect 504162 220170 504218 220226
rect 504038 220046 504094 220102
rect 504162 220046 504218 220102
rect 504038 219922 504094 219978
rect 504162 219922 504218 219978
rect 534758 220294 534814 220350
rect 534882 220294 534938 220350
rect 534758 220170 534814 220226
rect 534882 220170 534938 220226
rect 534758 220046 534814 220102
rect 534882 220046 534938 220102
rect 534758 219922 534814 219978
rect 534882 219922 534938 219978
rect 565478 220294 565534 220350
rect 565602 220294 565658 220350
rect 565478 220170 565534 220226
rect 565602 220170 565658 220226
rect 565478 220046 565534 220102
rect 565602 220046 565658 220102
rect 565478 219922 565534 219978
rect 565602 219922 565658 219978
rect 27878 208294 27934 208350
rect 28002 208294 28058 208350
rect 27878 208170 27934 208226
rect 28002 208170 28058 208226
rect 27878 208046 27934 208102
rect 28002 208046 28058 208102
rect 27878 207922 27934 207978
rect 28002 207922 28058 207978
rect 58598 208294 58654 208350
rect 58722 208294 58778 208350
rect 58598 208170 58654 208226
rect 58722 208170 58778 208226
rect 58598 208046 58654 208102
rect 58722 208046 58778 208102
rect 58598 207922 58654 207978
rect 58722 207922 58778 207978
rect 89318 208294 89374 208350
rect 89442 208294 89498 208350
rect 89318 208170 89374 208226
rect 89442 208170 89498 208226
rect 89318 208046 89374 208102
rect 89442 208046 89498 208102
rect 89318 207922 89374 207978
rect 89442 207922 89498 207978
rect 120038 208294 120094 208350
rect 120162 208294 120218 208350
rect 120038 208170 120094 208226
rect 120162 208170 120218 208226
rect 120038 208046 120094 208102
rect 120162 208046 120218 208102
rect 120038 207922 120094 207978
rect 120162 207922 120218 207978
rect 150758 208294 150814 208350
rect 150882 208294 150938 208350
rect 150758 208170 150814 208226
rect 150882 208170 150938 208226
rect 150758 208046 150814 208102
rect 150882 208046 150938 208102
rect 150758 207922 150814 207978
rect 150882 207922 150938 207978
rect 181478 208294 181534 208350
rect 181602 208294 181658 208350
rect 181478 208170 181534 208226
rect 181602 208170 181658 208226
rect 181478 208046 181534 208102
rect 181602 208046 181658 208102
rect 181478 207922 181534 207978
rect 181602 207922 181658 207978
rect 212198 208294 212254 208350
rect 212322 208294 212378 208350
rect 212198 208170 212254 208226
rect 212322 208170 212378 208226
rect 212198 208046 212254 208102
rect 212322 208046 212378 208102
rect 212198 207922 212254 207978
rect 212322 207922 212378 207978
rect 242918 208294 242974 208350
rect 243042 208294 243098 208350
rect 242918 208170 242974 208226
rect 243042 208170 243098 208226
rect 242918 208046 242974 208102
rect 243042 208046 243098 208102
rect 242918 207922 242974 207978
rect 243042 207922 243098 207978
rect 273638 208294 273694 208350
rect 273762 208294 273818 208350
rect 273638 208170 273694 208226
rect 273762 208170 273818 208226
rect 273638 208046 273694 208102
rect 273762 208046 273818 208102
rect 273638 207922 273694 207978
rect 273762 207922 273818 207978
rect 304358 208294 304414 208350
rect 304482 208294 304538 208350
rect 304358 208170 304414 208226
rect 304482 208170 304538 208226
rect 304358 208046 304414 208102
rect 304482 208046 304538 208102
rect 304358 207922 304414 207978
rect 304482 207922 304538 207978
rect 335078 208294 335134 208350
rect 335202 208294 335258 208350
rect 335078 208170 335134 208226
rect 335202 208170 335258 208226
rect 335078 208046 335134 208102
rect 335202 208046 335258 208102
rect 335078 207922 335134 207978
rect 335202 207922 335258 207978
rect 365798 208294 365854 208350
rect 365922 208294 365978 208350
rect 365798 208170 365854 208226
rect 365922 208170 365978 208226
rect 365798 208046 365854 208102
rect 365922 208046 365978 208102
rect 365798 207922 365854 207978
rect 365922 207922 365978 207978
rect 396518 208294 396574 208350
rect 396642 208294 396698 208350
rect 396518 208170 396574 208226
rect 396642 208170 396698 208226
rect 396518 208046 396574 208102
rect 396642 208046 396698 208102
rect 396518 207922 396574 207978
rect 396642 207922 396698 207978
rect 427238 208294 427294 208350
rect 427362 208294 427418 208350
rect 427238 208170 427294 208226
rect 427362 208170 427418 208226
rect 427238 208046 427294 208102
rect 427362 208046 427418 208102
rect 427238 207922 427294 207978
rect 427362 207922 427418 207978
rect 457958 208294 458014 208350
rect 458082 208294 458138 208350
rect 457958 208170 458014 208226
rect 458082 208170 458138 208226
rect 457958 208046 458014 208102
rect 458082 208046 458138 208102
rect 457958 207922 458014 207978
rect 458082 207922 458138 207978
rect 488678 208294 488734 208350
rect 488802 208294 488858 208350
rect 488678 208170 488734 208226
rect 488802 208170 488858 208226
rect 488678 208046 488734 208102
rect 488802 208046 488858 208102
rect 488678 207922 488734 207978
rect 488802 207922 488858 207978
rect 519398 208294 519454 208350
rect 519522 208294 519578 208350
rect 519398 208170 519454 208226
rect 519522 208170 519578 208226
rect 519398 208046 519454 208102
rect 519522 208046 519578 208102
rect 519398 207922 519454 207978
rect 519522 207922 519578 207978
rect 550118 208294 550174 208350
rect 550242 208294 550298 208350
rect 550118 208170 550174 208226
rect 550242 208170 550298 208226
rect 550118 208046 550174 208102
rect 550242 208046 550298 208102
rect 550118 207922 550174 207978
rect 550242 207922 550298 207978
rect 5514 202294 5570 202350
rect 5638 202294 5694 202350
rect 5762 202294 5818 202350
rect 5886 202294 5942 202350
rect 5514 202170 5570 202226
rect 5638 202170 5694 202226
rect 5762 202170 5818 202226
rect 5886 202170 5942 202226
rect 5514 202046 5570 202102
rect 5638 202046 5694 202102
rect 5762 202046 5818 202102
rect 5886 202046 5942 202102
rect 5514 201922 5570 201978
rect 5638 201922 5694 201978
rect 5762 201922 5818 201978
rect 5886 201922 5942 201978
rect -860 184294 -804 184350
rect -736 184294 -680 184350
rect -612 184294 -556 184350
rect -488 184294 -432 184350
rect -860 184170 -804 184226
rect -736 184170 -680 184226
rect -612 184170 -556 184226
rect -488 184170 -432 184226
rect -860 184046 -804 184102
rect -736 184046 -680 184102
rect -612 184046 -556 184102
rect -488 184046 -432 184102
rect -860 183922 -804 183978
rect -736 183922 -680 183978
rect -612 183922 -556 183978
rect -488 183922 -432 183978
rect 12518 202294 12574 202350
rect 12642 202294 12698 202350
rect 12518 202170 12574 202226
rect 12642 202170 12698 202226
rect 12518 202046 12574 202102
rect 12642 202046 12698 202102
rect 12518 201922 12574 201978
rect 12642 201922 12698 201978
rect 43238 202294 43294 202350
rect 43362 202294 43418 202350
rect 43238 202170 43294 202226
rect 43362 202170 43418 202226
rect 43238 202046 43294 202102
rect 43362 202046 43418 202102
rect 43238 201922 43294 201978
rect 43362 201922 43418 201978
rect 73958 202294 74014 202350
rect 74082 202294 74138 202350
rect 73958 202170 74014 202226
rect 74082 202170 74138 202226
rect 73958 202046 74014 202102
rect 74082 202046 74138 202102
rect 73958 201922 74014 201978
rect 74082 201922 74138 201978
rect 104678 202294 104734 202350
rect 104802 202294 104858 202350
rect 104678 202170 104734 202226
rect 104802 202170 104858 202226
rect 104678 202046 104734 202102
rect 104802 202046 104858 202102
rect 104678 201922 104734 201978
rect 104802 201922 104858 201978
rect 135398 202294 135454 202350
rect 135522 202294 135578 202350
rect 135398 202170 135454 202226
rect 135522 202170 135578 202226
rect 135398 202046 135454 202102
rect 135522 202046 135578 202102
rect 135398 201922 135454 201978
rect 135522 201922 135578 201978
rect 166118 202294 166174 202350
rect 166242 202294 166298 202350
rect 166118 202170 166174 202226
rect 166242 202170 166298 202226
rect 166118 202046 166174 202102
rect 166242 202046 166298 202102
rect 166118 201922 166174 201978
rect 166242 201922 166298 201978
rect 196838 202294 196894 202350
rect 196962 202294 197018 202350
rect 196838 202170 196894 202226
rect 196962 202170 197018 202226
rect 196838 202046 196894 202102
rect 196962 202046 197018 202102
rect 196838 201922 196894 201978
rect 196962 201922 197018 201978
rect 227558 202294 227614 202350
rect 227682 202294 227738 202350
rect 227558 202170 227614 202226
rect 227682 202170 227738 202226
rect 227558 202046 227614 202102
rect 227682 202046 227738 202102
rect 227558 201922 227614 201978
rect 227682 201922 227738 201978
rect 258278 202294 258334 202350
rect 258402 202294 258458 202350
rect 258278 202170 258334 202226
rect 258402 202170 258458 202226
rect 258278 202046 258334 202102
rect 258402 202046 258458 202102
rect 258278 201922 258334 201978
rect 258402 201922 258458 201978
rect 288998 202294 289054 202350
rect 289122 202294 289178 202350
rect 288998 202170 289054 202226
rect 289122 202170 289178 202226
rect 288998 202046 289054 202102
rect 289122 202046 289178 202102
rect 288998 201922 289054 201978
rect 289122 201922 289178 201978
rect 319718 202294 319774 202350
rect 319842 202294 319898 202350
rect 319718 202170 319774 202226
rect 319842 202170 319898 202226
rect 319718 202046 319774 202102
rect 319842 202046 319898 202102
rect 319718 201922 319774 201978
rect 319842 201922 319898 201978
rect 350438 202294 350494 202350
rect 350562 202294 350618 202350
rect 350438 202170 350494 202226
rect 350562 202170 350618 202226
rect 350438 202046 350494 202102
rect 350562 202046 350618 202102
rect 350438 201922 350494 201978
rect 350562 201922 350618 201978
rect 381158 202294 381214 202350
rect 381282 202294 381338 202350
rect 381158 202170 381214 202226
rect 381282 202170 381338 202226
rect 381158 202046 381214 202102
rect 381282 202046 381338 202102
rect 381158 201922 381214 201978
rect 381282 201922 381338 201978
rect 411878 202294 411934 202350
rect 412002 202294 412058 202350
rect 411878 202170 411934 202226
rect 412002 202170 412058 202226
rect 411878 202046 411934 202102
rect 412002 202046 412058 202102
rect 411878 201922 411934 201978
rect 412002 201922 412058 201978
rect 442598 202294 442654 202350
rect 442722 202294 442778 202350
rect 442598 202170 442654 202226
rect 442722 202170 442778 202226
rect 442598 202046 442654 202102
rect 442722 202046 442778 202102
rect 442598 201922 442654 201978
rect 442722 201922 442778 201978
rect 473318 202294 473374 202350
rect 473442 202294 473498 202350
rect 473318 202170 473374 202226
rect 473442 202170 473498 202226
rect 473318 202046 473374 202102
rect 473442 202046 473498 202102
rect 473318 201922 473374 201978
rect 473442 201922 473498 201978
rect 504038 202294 504094 202350
rect 504162 202294 504218 202350
rect 504038 202170 504094 202226
rect 504162 202170 504218 202226
rect 504038 202046 504094 202102
rect 504162 202046 504218 202102
rect 504038 201922 504094 201978
rect 504162 201922 504218 201978
rect 534758 202294 534814 202350
rect 534882 202294 534938 202350
rect 534758 202170 534814 202226
rect 534882 202170 534938 202226
rect 534758 202046 534814 202102
rect 534882 202046 534938 202102
rect 534758 201922 534814 201978
rect 534882 201922 534938 201978
rect 565478 202294 565534 202350
rect 565602 202294 565658 202350
rect 565478 202170 565534 202226
rect 565602 202170 565658 202226
rect 565478 202046 565534 202102
rect 565602 202046 565658 202102
rect 565478 201922 565534 201978
rect 565602 201922 565658 201978
rect 27878 190294 27934 190350
rect 28002 190294 28058 190350
rect 27878 190170 27934 190226
rect 28002 190170 28058 190226
rect 27878 190046 27934 190102
rect 28002 190046 28058 190102
rect 27878 189922 27934 189978
rect 28002 189922 28058 189978
rect 58598 190294 58654 190350
rect 58722 190294 58778 190350
rect 58598 190170 58654 190226
rect 58722 190170 58778 190226
rect 58598 190046 58654 190102
rect 58722 190046 58778 190102
rect 58598 189922 58654 189978
rect 58722 189922 58778 189978
rect 89318 190294 89374 190350
rect 89442 190294 89498 190350
rect 89318 190170 89374 190226
rect 89442 190170 89498 190226
rect 89318 190046 89374 190102
rect 89442 190046 89498 190102
rect 89318 189922 89374 189978
rect 89442 189922 89498 189978
rect 120038 190294 120094 190350
rect 120162 190294 120218 190350
rect 120038 190170 120094 190226
rect 120162 190170 120218 190226
rect 120038 190046 120094 190102
rect 120162 190046 120218 190102
rect 120038 189922 120094 189978
rect 120162 189922 120218 189978
rect 150758 190294 150814 190350
rect 150882 190294 150938 190350
rect 150758 190170 150814 190226
rect 150882 190170 150938 190226
rect 150758 190046 150814 190102
rect 150882 190046 150938 190102
rect 150758 189922 150814 189978
rect 150882 189922 150938 189978
rect 181478 190294 181534 190350
rect 181602 190294 181658 190350
rect 181478 190170 181534 190226
rect 181602 190170 181658 190226
rect 181478 190046 181534 190102
rect 181602 190046 181658 190102
rect 181478 189922 181534 189978
rect 181602 189922 181658 189978
rect 212198 190294 212254 190350
rect 212322 190294 212378 190350
rect 212198 190170 212254 190226
rect 212322 190170 212378 190226
rect 212198 190046 212254 190102
rect 212322 190046 212378 190102
rect 212198 189922 212254 189978
rect 212322 189922 212378 189978
rect 242918 190294 242974 190350
rect 243042 190294 243098 190350
rect 242918 190170 242974 190226
rect 243042 190170 243098 190226
rect 242918 190046 242974 190102
rect 243042 190046 243098 190102
rect 242918 189922 242974 189978
rect 243042 189922 243098 189978
rect 273638 190294 273694 190350
rect 273762 190294 273818 190350
rect 273638 190170 273694 190226
rect 273762 190170 273818 190226
rect 273638 190046 273694 190102
rect 273762 190046 273818 190102
rect 273638 189922 273694 189978
rect 273762 189922 273818 189978
rect 304358 190294 304414 190350
rect 304482 190294 304538 190350
rect 304358 190170 304414 190226
rect 304482 190170 304538 190226
rect 304358 190046 304414 190102
rect 304482 190046 304538 190102
rect 304358 189922 304414 189978
rect 304482 189922 304538 189978
rect 335078 190294 335134 190350
rect 335202 190294 335258 190350
rect 335078 190170 335134 190226
rect 335202 190170 335258 190226
rect 335078 190046 335134 190102
rect 335202 190046 335258 190102
rect 335078 189922 335134 189978
rect 335202 189922 335258 189978
rect 365798 190294 365854 190350
rect 365922 190294 365978 190350
rect 365798 190170 365854 190226
rect 365922 190170 365978 190226
rect 365798 190046 365854 190102
rect 365922 190046 365978 190102
rect 365798 189922 365854 189978
rect 365922 189922 365978 189978
rect 396518 190294 396574 190350
rect 396642 190294 396698 190350
rect 396518 190170 396574 190226
rect 396642 190170 396698 190226
rect 396518 190046 396574 190102
rect 396642 190046 396698 190102
rect 396518 189922 396574 189978
rect 396642 189922 396698 189978
rect 427238 190294 427294 190350
rect 427362 190294 427418 190350
rect 427238 190170 427294 190226
rect 427362 190170 427418 190226
rect 427238 190046 427294 190102
rect 427362 190046 427418 190102
rect 427238 189922 427294 189978
rect 427362 189922 427418 189978
rect 457958 190294 458014 190350
rect 458082 190294 458138 190350
rect 457958 190170 458014 190226
rect 458082 190170 458138 190226
rect 457958 190046 458014 190102
rect 458082 190046 458138 190102
rect 457958 189922 458014 189978
rect 458082 189922 458138 189978
rect 488678 190294 488734 190350
rect 488802 190294 488858 190350
rect 488678 190170 488734 190226
rect 488802 190170 488858 190226
rect 488678 190046 488734 190102
rect 488802 190046 488858 190102
rect 488678 189922 488734 189978
rect 488802 189922 488858 189978
rect 519398 190294 519454 190350
rect 519522 190294 519578 190350
rect 519398 190170 519454 190226
rect 519522 190170 519578 190226
rect 519398 190046 519454 190102
rect 519522 190046 519578 190102
rect 519398 189922 519454 189978
rect 519522 189922 519578 189978
rect 550118 190294 550174 190350
rect 550242 190294 550298 190350
rect 550118 190170 550174 190226
rect 550242 190170 550298 190226
rect 550118 190046 550174 190102
rect 550242 190046 550298 190102
rect 550118 189922 550174 189978
rect 550242 189922 550298 189978
rect 5514 184294 5570 184350
rect 5638 184294 5694 184350
rect 5762 184294 5818 184350
rect 5886 184294 5942 184350
rect 5514 184170 5570 184226
rect 5638 184170 5694 184226
rect 5762 184170 5818 184226
rect 5886 184170 5942 184226
rect 5514 184046 5570 184102
rect 5638 184046 5694 184102
rect 5762 184046 5818 184102
rect 5886 184046 5942 184102
rect 5514 183922 5570 183978
rect 5638 183922 5694 183978
rect 5762 183922 5818 183978
rect 5886 183922 5942 183978
rect -860 166294 -804 166350
rect -736 166294 -680 166350
rect -612 166294 -556 166350
rect -488 166294 -432 166350
rect -860 166170 -804 166226
rect -736 166170 -680 166226
rect -612 166170 -556 166226
rect -488 166170 -432 166226
rect -860 166046 -804 166102
rect -736 166046 -680 166102
rect -612 166046 -556 166102
rect -488 166046 -432 166102
rect -860 165922 -804 165978
rect -736 165922 -680 165978
rect -612 165922 -556 165978
rect -488 165922 -432 165978
rect 12518 184294 12574 184350
rect 12642 184294 12698 184350
rect 12518 184170 12574 184226
rect 12642 184170 12698 184226
rect 12518 184046 12574 184102
rect 12642 184046 12698 184102
rect 12518 183922 12574 183978
rect 12642 183922 12698 183978
rect 43238 184294 43294 184350
rect 43362 184294 43418 184350
rect 43238 184170 43294 184226
rect 43362 184170 43418 184226
rect 43238 184046 43294 184102
rect 43362 184046 43418 184102
rect 43238 183922 43294 183978
rect 43362 183922 43418 183978
rect 73958 184294 74014 184350
rect 74082 184294 74138 184350
rect 73958 184170 74014 184226
rect 74082 184170 74138 184226
rect 73958 184046 74014 184102
rect 74082 184046 74138 184102
rect 73958 183922 74014 183978
rect 74082 183922 74138 183978
rect 104678 184294 104734 184350
rect 104802 184294 104858 184350
rect 104678 184170 104734 184226
rect 104802 184170 104858 184226
rect 104678 184046 104734 184102
rect 104802 184046 104858 184102
rect 104678 183922 104734 183978
rect 104802 183922 104858 183978
rect 135398 184294 135454 184350
rect 135522 184294 135578 184350
rect 135398 184170 135454 184226
rect 135522 184170 135578 184226
rect 135398 184046 135454 184102
rect 135522 184046 135578 184102
rect 135398 183922 135454 183978
rect 135522 183922 135578 183978
rect 166118 184294 166174 184350
rect 166242 184294 166298 184350
rect 166118 184170 166174 184226
rect 166242 184170 166298 184226
rect 166118 184046 166174 184102
rect 166242 184046 166298 184102
rect 166118 183922 166174 183978
rect 166242 183922 166298 183978
rect 196838 184294 196894 184350
rect 196962 184294 197018 184350
rect 196838 184170 196894 184226
rect 196962 184170 197018 184226
rect 196838 184046 196894 184102
rect 196962 184046 197018 184102
rect 196838 183922 196894 183978
rect 196962 183922 197018 183978
rect 227558 184294 227614 184350
rect 227682 184294 227738 184350
rect 227558 184170 227614 184226
rect 227682 184170 227738 184226
rect 227558 184046 227614 184102
rect 227682 184046 227738 184102
rect 227558 183922 227614 183978
rect 227682 183922 227738 183978
rect 258278 184294 258334 184350
rect 258402 184294 258458 184350
rect 258278 184170 258334 184226
rect 258402 184170 258458 184226
rect 258278 184046 258334 184102
rect 258402 184046 258458 184102
rect 258278 183922 258334 183978
rect 258402 183922 258458 183978
rect 288998 184294 289054 184350
rect 289122 184294 289178 184350
rect 288998 184170 289054 184226
rect 289122 184170 289178 184226
rect 288998 184046 289054 184102
rect 289122 184046 289178 184102
rect 288998 183922 289054 183978
rect 289122 183922 289178 183978
rect 319718 184294 319774 184350
rect 319842 184294 319898 184350
rect 319718 184170 319774 184226
rect 319842 184170 319898 184226
rect 319718 184046 319774 184102
rect 319842 184046 319898 184102
rect 319718 183922 319774 183978
rect 319842 183922 319898 183978
rect 350438 184294 350494 184350
rect 350562 184294 350618 184350
rect 350438 184170 350494 184226
rect 350562 184170 350618 184226
rect 350438 184046 350494 184102
rect 350562 184046 350618 184102
rect 350438 183922 350494 183978
rect 350562 183922 350618 183978
rect 381158 184294 381214 184350
rect 381282 184294 381338 184350
rect 381158 184170 381214 184226
rect 381282 184170 381338 184226
rect 381158 184046 381214 184102
rect 381282 184046 381338 184102
rect 381158 183922 381214 183978
rect 381282 183922 381338 183978
rect 411878 184294 411934 184350
rect 412002 184294 412058 184350
rect 411878 184170 411934 184226
rect 412002 184170 412058 184226
rect 411878 184046 411934 184102
rect 412002 184046 412058 184102
rect 411878 183922 411934 183978
rect 412002 183922 412058 183978
rect 442598 184294 442654 184350
rect 442722 184294 442778 184350
rect 442598 184170 442654 184226
rect 442722 184170 442778 184226
rect 442598 184046 442654 184102
rect 442722 184046 442778 184102
rect 442598 183922 442654 183978
rect 442722 183922 442778 183978
rect 473318 184294 473374 184350
rect 473442 184294 473498 184350
rect 473318 184170 473374 184226
rect 473442 184170 473498 184226
rect 473318 184046 473374 184102
rect 473442 184046 473498 184102
rect 473318 183922 473374 183978
rect 473442 183922 473498 183978
rect 504038 184294 504094 184350
rect 504162 184294 504218 184350
rect 504038 184170 504094 184226
rect 504162 184170 504218 184226
rect 504038 184046 504094 184102
rect 504162 184046 504218 184102
rect 504038 183922 504094 183978
rect 504162 183922 504218 183978
rect 534758 184294 534814 184350
rect 534882 184294 534938 184350
rect 534758 184170 534814 184226
rect 534882 184170 534938 184226
rect 534758 184046 534814 184102
rect 534882 184046 534938 184102
rect 534758 183922 534814 183978
rect 534882 183922 534938 183978
rect 565478 184294 565534 184350
rect 565602 184294 565658 184350
rect 565478 184170 565534 184226
rect 565602 184170 565658 184226
rect 565478 184046 565534 184102
rect 565602 184046 565658 184102
rect 565478 183922 565534 183978
rect 565602 183922 565658 183978
rect 592914 280294 592970 280350
rect 593038 280294 593094 280350
rect 593162 280294 593218 280350
rect 593286 280294 593342 280350
rect 592914 280170 592970 280226
rect 593038 280170 593094 280226
rect 593162 280170 593218 280226
rect 593286 280170 593342 280226
rect 592914 280046 592970 280102
rect 593038 280046 593094 280102
rect 593162 280046 593218 280102
rect 593286 280046 593342 280102
rect 592914 279922 592970 279978
rect 593038 279922 593094 279978
rect 593162 279922 593218 279978
rect 593286 279922 593342 279978
rect 589194 256294 589250 256350
rect 589318 256294 589374 256350
rect 589442 256294 589498 256350
rect 589566 256294 589622 256350
rect 589194 256170 589250 256226
rect 589318 256170 589374 256226
rect 589442 256170 589498 256226
rect 589566 256170 589622 256226
rect 589194 256046 589250 256102
rect 589318 256046 589374 256102
rect 589442 256046 589498 256102
rect 589566 256046 589622 256102
rect 589194 255922 589250 255978
rect 589318 255922 589374 255978
rect 589442 255922 589498 255978
rect 589566 255922 589622 255978
rect 592914 262294 592970 262350
rect 593038 262294 593094 262350
rect 593162 262294 593218 262350
rect 593286 262294 593342 262350
rect 592914 262170 592970 262226
rect 593038 262170 593094 262226
rect 593162 262170 593218 262226
rect 593286 262170 593342 262226
rect 592914 262046 592970 262102
rect 593038 262046 593094 262102
rect 593162 262046 593218 262102
rect 593286 262046 593342 262102
rect 592914 261922 592970 261978
rect 593038 261922 593094 261978
rect 593162 261922 593218 261978
rect 593286 261922 593342 261978
rect 589194 238294 589250 238350
rect 589318 238294 589374 238350
rect 589442 238294 589498 238350
rect 589566 238294 589622 238350
rect 589194 238170 589250 238226
rect 589318 238170 589374 238226
rect 589442 238170 589498 238226
rect 589566 238170 589622 238226
rect 589194 238046 589250 238102
rect 589318 238046 589374 238102
rect 589442 238046 589498 238102
rect 589566 238046 589622 238102
rect 589194 237922 589250 237978
rect 589318 237922 589374 237978
rect 589442 237922 589498 237978
rect 589566 237922 589622 237978
rect 589194 220294 589250 220350
rect 589318 220294 589374 220350
rect 589442 220294 589498 220350
rect 589566 220294 589622 220350
rect 589194 220170 589250 220226
rect 589318 220170 589374 220226
rect 589442 220170 589498 220226
rect 589566 220170 589622 220226
rect 589194 220046 589250 220102
rect 589318 220046 589374 220102
rect 589442 220046 589498 220102
rect 589566 220046 589622 220102
rect 589194 219922 589250 219978
rect 589318 219922 589374 219978
rect 589442 219922 589498 219978
rect 589566 219922 589622 219978
rect 592914 244294 592970 244350
rect 593038 244294 593094 244350
rect 593162 244294 593218 244350
rect 593286 244294 593342 244350
rect 592914 244170 592970 244226
rect 593038 244170 593094 244226
rect 593162 244170 593218 244226
rect 593286 244170 593342 244226
rect 592914 244046 592970 244102
rect 593038 244046 593094 244102
rect 593162 244046 593218 244102
rect 593286 244046 593342 244102
rect 592914 243922 592970 243978
rect 593038 243922 593094 243978
rect 593162 243922 593218 243978
rect 593286 243922 593342 243978
rect 592914 226294 592970 226350
rect 593038 226294 593094 226350
rect 593162 226294 593218 226350
rect 593286 226294 593342 226350
rect 592914 226170 592970 226226
rect 593038 226170 593094 226226
rect 593162 226170 593218 226226
rect 593286 226170 593342 226226
rect 592914 226046 592970 226102
rect 593038 226046 593094 226102
rect 593162 226046 593218 226102
rect 593286 226046 593342 226102
rect 592914 225922 592970 225978
rect 593038 225922 593094 225978
rect 593162 225922 593218 225978
rect 593286 225922 593342 225978
rect 589194 202294 589250 202350
rect 589318 202294 589374 202350
rect 589442 202294 589498 202350
rect 589566 202294 589622 202350
rect 589194 202170 589250 202226
rect 589318 202170 589374 202226
rect 589442 202170 589498 202226
rect 589566 202170 589622 202226
rect 589194 202046 589250 202102
rect 589318 202046 589374 202102
rect 589442 202046 589498 202102
rect 589566 202046 589622 202102
rect 589194 201922 589250 201978
rect 589318 201922 589374 201978
rect 589442 201922 589498 201978
rect 589566 201922 589622 201978
rect 27878 172294 27934 172350
rect 28002 172294 28058 172350
rect 27878 172170 27934 172226
rect 28002 172170 28058 172226
rect 27878 172046 27934 172102
rect 28002 172046 28058 172102
rect 27878 171922 27934 171978
rect 28002 171922 28058 171978
rect 58598 172294 58654 172350
rect 58722 172294 58778 172350
rect 58598 172170 58654 172226
rect 58722 172170 58778 172226
rect 58598 172046 58654 172102
rect 58722 172046 58778 172102
rect 58598 171922 58654 171978
rect 58722 171922 58778 171978
rect 89318 172294 89374 172350
rect 89442 172294 89498 172350
rect 89318 172170 89374 172226
rect 89442 172170 89498 172226
rect 89318 172046 89374 172102
rect 89442 172046 89498 172102
rect 89318 171922 89374 171978
rect 89442 171922 89498 171978
rect 120038 172294 120094 172350
rect 120162 172294 120218 172350
rect 120038 172170 120094 172226
rect 120162 172170 120218 172226
rect 120038 172046 120094 172102
rect 120162 172046 120218 172102
rect 120038 171922 120094 171978
rect 120162 171922 120218 171978
rect 150758 172294 150814 172350
rect 150882 172294 150938 172350
rect 150758 172170 150814 172226
rect 150882 172170 150938 172226
rect 150758 172046 150814 172102
rect 150882 172046 150938 172102
rect 150758 171922 150814 171978
rect 150882 171922 150938 171978
rect 181478 172294 181534 172350
rect 181602 172294 181658 172350
rect 181478 172170 181534 172226
rect 181602 172170 181658 172226
rect 181478 172046 181534 172102
rect 181602 172046 181658 172102
rect 181478 171922 181534 171978
rect 181602 171922 181658 171978
rect 212198 172294 212254 172350
rect 212322 172294 212378 172350
rect 212198 172170 212254 172226
rect 212322 172170 212378 172226
rect 212198 172046 212254 172102
rect 212322 172046 212378 172102
rect 212198 171922 212254 171978
rect 212322 171922 212378 171978
rect 242918 172294 242974 172350
rect 243042 172294 243098 172350
rect 242918 172170 242974 172226
rect 243042 172170 243098 172226
rect 242918 172046 242974 172102
rect 243042 172046 243098 172102
rect 242918 171922 242974 171978
rect 243042 171922 243098 171978
rect 273638 172294 273694 172350
rect 273762 172294 273818 172350
rect 273638 172170 273694 172226
rect 273762 172170 273818 172226
rect 273638 172046 273694 172102
rect 273762 172046 273818 172102
rect 273638 171922 273694 171978
rect 273762 171922 273818 171978
rect 304358 172294 304414 172350
rect 304482 172294 304538 172350
rect 304358 172170 304414 172226
rect 304482 172170 304538 172226
rect 304358 172046 304414 172102
rect 304482 172046 304538 172102
rect 304358 171922 304414 171978
rect 304482 171922 304538 171978
rect 335078 172294 335134 172350
rect 335202 172294 335258 172350
rect 335078 172170 335134 172226
rect 335202 172170 335258 172226
rect 335078 172046 335134 172102
rect 335202 172046 335258 172102
rect 335078 171922 335134 171978
rect 335202 171922 335258 171978
rect 365798 172294 365854 172350
rect 365922 172294 365978 172350
rect 365798 172170 365854 172226
rect 365922 172170 365978 172226
rect 365798 172046 365854 172102
rect 365922 172046 365978 172102
rect 365798 171922 365854 171978
rect 365922 171922 365978 171978
rect 396518 172294 396574 172350
rect 396642 172294 396698 172350
rect 396518 172170 396574 172226
rect 396642 172170 396698 172226
rect 396518 172046 396574 172102
rect 396642 172046 396698 172102
rect 396518 171922 396574 171978
rect 396642 171922 396698 171978
rect 427238 172294 427294 172350
rect 427362 172294 427418 172350
rect 427238 172170 427294 172226
rect 427362 172170 427418 172226
rect 427238 172046 427294 172102
rect 427362 172046 427418 172102
rect 427238 171922 427294 171978
rect 427362 171922 427418 171978
rect 457958 172294 458014 172350
rect 458082 172294 458138 172350
rect 457958 172170 458014 172226
rect 458082 172170 458138 172226
rect 457958 172046 458014 172102
rect 458082 172046 458138 172102
rect 457958 171922 458014 171978
rect 458082 171922 458138 171978
rect 488678 172294 488734 172350
rect 488802 172294 488858 172350
rect 488678 172170 488734 172226
rect 488802 172170 488858 172226
rect 488678 172046 488734 172102
rect 488802 172046 488858 172102
rect 488678 171922 488734 171978
rect 488802 171922 488858 171978
rect 519398 172294 519454 172350
rect 519522 172294 519578 172350
rect 519398 172170 519454 172226
rect 519522 172170 519578 172226
rect 519398 172046 519454 172102
rect 519522 172046 519578 172102
rect 519398 171922 519454 171978
rect 519522 171922 519578 171978
rect 550118 172294 550174 172350
rect 550242 172294 550298 172350
rect 550118 172170 550174 172226
rect 550242 172170 550298 172226
rect 550118 172046 550174 172102
rect 550242 172046 550298 172102
rect 550118 171922 550174 171978
rect 550242 171922 550298 171978
rect 589194 184294 589250 184350
rect 589318 184294 589374 184350
rect 589442 184294 589498 184350
rect 589566 184294 589622 184350
rect 589194 184170 589250 184226
rect 589318 184170 589374 184226
rect 589442 184170 589498 184226
rect 589566 184170 589622 184226
rect 589194 184046 589250 184102
rect 589318 184046 589374 184102
rect 589442 184046 589498 184102
rect 589566 184046 589622 184102
rect 589194 183922 589250 183978
rect 589318 183922 589374 183978
rect 589442 183922 589498 183978
rect 589566 183922 589622 183978
rect 5514 166294 5570 166350
rect 5638 166294 5694 166350
rect 5762 166294 5818 166350
rect 5886 166294 5942 166350
rect 5514 166170 5570 166226
rect 5638 166170 5694 166226
rect 5762 166170 5818 166226
rect 5886 166170 5942 166226
rect 5514 166046 5570 166102
rect 5638 166046 5694 166102
rect 5762 166046 5818 166102
rect 5886 166046 5942 166102
rect 5514 165922 5570 165978
rect 5638 165922 5694 165978
rect 5762 165922 5818 165978
rect 5886 165922 5942 165978
rect -860 148294 -804 148350
rect -736 148294 -680 148350
rect -612 148294 -556 148350
rect -488 148294 -432 148350
rect -860 148170 -804 148226
rect -736 148170 -680 148226
rect -612 148170 -556 148226
rect -488 148170 -432 148226
rect -860 148046 -804 148102
rect -736 148046 -680 148102
rect -612 148046 -556 148102
rect -488 148046 -432 148102
rect -860 147922 -804 147978
rect -736 147922 -680 147978
rect -612 147922 -556 147978
rect -488 147922 -432 147978
rect 12518 166294 12574 166350
rect 12642 166294 12698 166350
rect 12518 166170 12574 166226
rect 12642 166170 12698 166226
rect 12518 166046 12574 166102
rect 12642 166046 12698 166102
rect 12518 165922 12574 165978
rect 12642 165922 12698 165978
rect 43238 166294 43294 166350
rect 43362 166294 43418 166350
rect 43238 166170 43294 166226
rect 43362 166170 43418 166226
rect 43238 166046 43294 166102
rect 43362 166046 43418 166102
rect 43238 165922 43294 165978
rect 43362 165922 43418 165978
rect 73958 166294 74014 166350
rect 74082 166294 74138 166350
rect 73958 166170 74014 166226
rect 74082 166170 74138 166226
rect 73958 166046 74014 166102
rect 74082 166046 74138 166102
rect 73958 165922 74014 165978
rect 74082 165922 74138 165978
rect 104678 166294 104734 166350
rect 104802 166294 104858 166350
rect 104678 166170 104734 166226
rect 104802 166170 104858 166226
rect 104678 166046 104734 166102
rect 104802 166046 104858 166102
rect 104678 165922 104734 165978
rect 104802 165922 104858 165978
rect 135398 166294 135454 166350
rect 135522 166294 135578 166350
rect 135398 166170 135454 166226
rect 135522 166170 135578 166226
rect 135398 166046 135454 166102
rect 135522 166046 135578 166102
rect 135398 165922 135454 165978
rect 135522 165922 135578 165978
rect 166118 166294 166174 166350
rect 166242 166294 166298 166350
rect 166118 166170 166174 166226
rect 166242 166170 166298 166226
rect 166118 166046 166174 166102
rect 166242 166046 166298 166102
rect 166118 165922 166174 165978
rect 166242 165922 166298 165978
rect 196838 166294 196894 166350
rect 196962 166294 197018 166350
rect 196838 166170 196894 166226
rect 196962 166170 197018 166226
rect 196838 166046 196894 166102
rect 196962 166046 197018 166102
rect 196838 165922 196894 165978
rect 196962 165922 197018 165978
rect 227558 166294 227614 166350
rect 227682 166294 227738 166350
rect 227558 166170 227614 166226
rect 227682 166170 227738 166226
rect 227558 166046 227614 166102
rect 227682 166046 227738 166102
rect 227558 165922 227614 165978
rect 227682 165922 227738 165978
rect 258278 166294 258334 166350
rect 258402 166294 258458 166350
rect 258278 166170 258334 166226
rect 258402 166170 258458 166226
rect 258278 166046 258334 166102
rect 258402 166046 258458 166102
rect 258278 165922 258334 165978
rect 258402 165922 258458 165978
rect 288998 166294 289054 166350
rect 289122 166294 289178 166350
rect 288998 166170 289054 166226
rect 289122 166170 289178 166226
rect 288998 166046 289054 166102
rect 289122 166046 289178 166102
rect 288998 165922 289054 165978
rect 289122 165922 289178 165978
rect 319718 166294 319774 166350
rect 319842 166294 319898 166350
rect 319718 166170 319774 166226
rect 319842 166170 319898 166226
rect 319718 166046 319774 166102
rect 319842 166046 319898 166102
rect 319718 165922 319774 165978
rect 319842 165922 319898 165978
rect 350438 166294 350494 166350
rect 350562 166294 350618 166350
rect 350438 166170 350494 166226
rect 350562 166170 350618 166226
rect 350438 166046 350494 166102
rect 350562 166046 350618 166102
rect 350438 165922 350494 165978
rect 350562 165922 350618 165978
rect 381158 166294 381214 166350
rect 381282 166294 381338 166350
rect 381158 166170 381214 166226
rect 381282 166170 381338 166226
rect 381158 166046 381214 166102
rect 381282 166046 381338 166102
rect 381158 165922 381214 165978
rect 381282 165922 381338 165978
rect 411878 166294 411934 166350
rect 412002 166294 412058 166350
rect 411878 166170 411934 166226
rect 412002 166170 412058 166226
rect 411878 166046 411934 166102
rect 412002 166046 412058 166102
rect 411878 165922 411934 165978
rect 412002 165922 412058 165978
rect 442598 166294 442654 166350
rect 442722 166294 442778 166350
rect 442598 166170 442654 166226
rect 442722 166170 442778 166226
rect 442598 166046 442654 166102
rect 442722 166046 442778 166102
rect 442598 165922 442654 165978
rect 442722 165922 442778 165978
rect 473318 166294 473374 166350
rect 473442 166294 473498 166350
rect 473318 166170 473374 166226
rect 473442 166170 473498 166226
rect 473318 166046 473374 166102
rect 473442 166046 473498 166102
rect 473318 165922 473374 165978
rect 473442 165922 473498 165978
rect 504038 166294 504094 166350
rect 504162 166294 504218 166350
rect 504038 166170 504094 166226
rect 504162 166170 504218 166226
rect 504038 166046 504094 166102
rect 504162 166046 504218 166102
rect 504038 165922 504094 165978
rect 504162 165922 504218 165978
rect 534758 166294 534814 166350
rect 534882 166294 534938 166350
rect 534758 166170 534814 166226
rect 534882 166170 534938 166226
rect 534758 166046 534814 166102
rect 534882 166046 534938 166102
rect 534758 165922 534814 165978
rect 534882 165922 534938 165978
rect 565478 166294 565534 166350
rect 565602 166294 565658 166350
rect 565478 166170 565534 166226
rect 565602 166170 565658 166226
rect 565478 166046 565534 166102
rect 565602 166046 565658 166102
rect 565478 165922 565534 165978
rect 565602 165922 565658 165978
rect 5514 148294 5570 148350
rect 5638 148294 5694 148350
rect 5762 148294 5818 148350
rect 5886 148294 5942 148350
rect 5514 148170 5570 148226
rect 5638 148170 5694 148226
rect 5762 148170 5818 148226
rect 5886 148170 5942 148226
rect 5514 148046 5570 148102
rect 5638 148046 5694 148102
rect 5762 148046 5818 148102
rect 5886 148046 5942 148102
rect 5514 147922 5570 147978
rect 5638 147922 5694 147978
rect 5762 147922 5818 147978
rect 5886 147922 5942 147978
rect -860 130294 -804 130350
rect -736 130294 -680 130350
rect -612 130294 -556 130350
rect -488 130294 -432 130350
rect -860 130170 -804 130226
rect -736 130170 -680 130226
rect -612 130170 -556 130226
rect -488 130170 -432 130226
rect -860 130046 -804 130102
rect -736 130046 -680 130102
rect -612 130046 -556 130102
rect -488 130046 -432 130102
rect -860 129922 -804 129978
rect -736 129922 -680 129978
rect -612 129922 -556 129978
rect -488 129922 -432 129978
rect 27878 154294 27934 154350
rect 28002 154294 28058 154350
rect 27878 154170 27934 154226
rect 28002 154170 28058 154226
rect 27878 154046 27934 154102
rect 28002 154046 28058 154102
rect 27878 153922 27934 153978
rect 28002 153922 28058 153978
rect 58598 154294 58654 154350
rect 58722 154294 58778 154350
rect 58598 154170 58654 154226
rect 58722 154170 58778 154226
rect 58598 154046 58654 154102
rect 58722 154046 58778 154102
rect 58598 153922 58654 153978
rect 58722 153922 58778 153978
rect 89318 154294 89374 154350
rect 89442 154294 89498 154350
rect 89318 154170 89374 154226
rect 89442 154170 89498 154226
rect 89318 154046 89374 154102
rect 89442 154046 89498 154102
rect 89318 153922 89374 153978
rect 89442 153922 89498 153978
rect 120038 154294 120094 154350
rect 120162 154294 120218 154350
rect 120038 154170 120094 154226
rect 120162 154170 120218 154226
rect 120038 154046 120094 154102
rect 120162 154046 120218 154102
rect 120038 153922 120094 153978
rect 120162 153922 120218 153978
rect 150758 154294 150814 154350
rect 150882 154294 150938 154350
rect 150758 154170 150814 154226
rect 150882 154170 150938 154226
rect 150758 154046 150814 154102
rect 150882 154046 150938 154102
rect 150758 153922 150814 153978
rect 150882 153922 150938 153978
rect 181478 154294 181534 154350
rect 181602 154294 181658 154350
rect 181478 154170 181534 154226
rect 181602 154170 181658 154226
rect 181478 154046 181534 154102
rect 181602 154046 181658 154102
rect 181478 153922 181534 153978
rect 181602 153922 181658 153978
rect 212198 154294 212254 154350
rect 212322 154294 212378 154350
rect 212198 154170 212254 154226
rect 212322 154170 212378 154226
rect 212198 154046 212254 154102
rect 212322 154046 212378 154102
rect 212198 153922 212254 153978
rect 212322 153922 212378 153978
rect 242918 154294 242974 154350
rect 243042 154294 243098 154350
rect 242918 154170 242974 154226
rect 243042 154170 243098 154226
rect 242918 154046 242974 154102
rect 243042 154046 243098 154102
rect 242918 153922 242974 153978
rect 243042 153922 243098 153978
rect 273638 154294 273694 154350
rect 273762 154294 273818 154350
rect 273638 154170 273694 154226
rect 273762 154170 273818 154226
rect 273638 154046 273694 154102
rect 273762 154046 273818 154102
rect 273638 153922 273694 153978
rect 273762 153922 273818 153978
rect 304358 154294 304414 154350
rect 304482 154294 304538 154350
rect 304358 154170 304414 154226
rect 304482 154170 304538 154226
rect 304358 154046 304414 154102
rect 304482 154046 304538 154102
rect 304358 153922 304414 153978
rect 304482 153922 304538 153978
rect 335078 154294 335134 154350
rect 335202 154294 335258 154350
rect 335078 154170 335134 154226
rect 335202 154170 335258 154226
rect 335078 154046 335134 154102
rect 335202 154046 335258 154102
rect 335078 153922 335134 153978
rect 335202 153922 335258 153978
rect 365798 154294 365854 154350
rect 365922 154294 365978 154350
rect 365798 154170 365854 154226
rect 365922 154170 365978 154226
rect 365798 154046 365854 154102
rect 365922 154046 365978 154102
rect 365798 153922 365854 153978
rect 365922 153922 365978 153978
rect 396518 154294 396574 154350
rect 396642 154294 396698 154350
rect 396518 154170 396574 154226
rect 396642 154170 396698 154226
rect 396518 154046 396574 154102
rect 396642 154046 396698 154102
rect 396518 153922 396574 153978
rect 396642 153922 396698 153978
rect 427238 154294 427294 154350
rect 427362 154294 427418 154350
rect 427238 154170 427294 154226
rect 427362 154170 427418 154226
rect 427238 154046 427294 154102
rect 427362 154046 427418 154102
rect 427238 153922 427294 153978
rect 427362 153922 427418 153978
rect 457958 154294 458014 154350
rect 458082 154294 458138 154350
rect 457958 154170 458014 154226
rect 458082 154170 458138 154226
rect 457958 154046 458014 154102
rect 458082 154046 458138 154102
rect 457958 153922 458014 153978
rect 458082 153922 458138 153978
rect 488678 154294 488734 154350
rect 488802 154294 488858 154350
rect 488678 154170 488734 154226
rect 488802 154170 488858 154226
rect 488678 154046 488734 154102
rect 488802 154046 488858 154102
rect 488678 153922 488734 153978
rect 488802 153922 488858 153978
rect 519398 154294 519454 154350
rect 519522 154294 519578 154350
rect 519398 154170 519454 154226
rect 519522 154170 519578 154226
rect 519398 154046 519454 154102
rect 519522 154046 519578 154102
rect 519398 153922 519454 153978
rect 519522 153922 519578 153978
rect 550118 154294 550174 154350
rect 550242 154294 550298 154350
rect 550118 154170 550174 154226
rect 550242 154170 550298 154226
rect 550118 154046 550174 154102
rect 550242 154046 550298 154102
rect 550118 153922 550174 153978
rect 550242 153922 550298 153978
rect 12518 148294 12574 148350
rect 12642 148294 12698 148350
rect 12518 148170 12574 148226
rect 12642 148170 12698 148226
rect 12518 148046 12574 148102
rect 12642 148046 12698 148102
rect 12518 147922 12574 147978
rect 12642 147922 12698 147978
rect 43238 148294 43294 148350
rect 43362 148294 43418 148350
rect 43238 148170 43294 148226
rect 43362 148170 43418 148226
rect 43238 148046 43294 148102
rect 43362 148046 43418 148102
rect 43238 147922 43294 147978
rect 43362 147922 43418 147978
rect 73958 148294 74014 148350
rect 74082 148294 74138 148350
rect 73958 148170 74014 148226
rect 74082 148170 74138 148226
rect 73958 148046 74014 148102
rect 74082 148046 74138 148102
rect 73958 147922 74014 147978
rect 74082 147922 74138 147978
rect 104678 148294 104734 148350
rect 104802 148294 104858 148350
rect 104678 148170 104734 148226
rect 104802 148170 104858 148226
rect 104678 148046 104734 148102
rect 104802 148046 104858 148102
rect 104678 147922 104734 147978
rect 104802 147922 104858 147978
rect 135398 148294 135454 148350
rect 135522 148294 135578 148350
rect 135398 148170 135454 148226
rect 135522 148170 135578 148226
rect 135398 148046 135454 148102
rect 135522 148046 135578 148102
rect 135398 147922 135454 147978
rect 135522 147922 135578 147978
rect 166118 148294 166174 148350
rect 166242 148294 166298 148350
rect 166118 148170 166174 148226
rect 166242 148170 166298 148226
rect 166118 148046 166174 148102
rect 166242 148046 166298 148102
rect 166118 147922 166174 147978
rect 166242 147922 166298 147978
rect 196838 148294 196894 148350
rect 196962 148294 197018 148350
rect 196838 148170 196894 148226
rect 196962 148170 197018 148226
rect 196838 148046 196894 148102
rect 196962 148046 197018 148102
rect 196838 147922 196894 147978
rect 196962 147922 197018 147978
rect 227558 148294 227614 148350
rect 227682 148294 227738 148350
rect 227558 148170 227614 148226
rect 227682 148170 227738 148226
rect 227558 148046 227614 148102
rect 227682 148046 227738 148102
rect 227558 147922 227614 147978
rect 227682 147922 227738 147978
rect 258278 148294 258334 148350
rect 258402 148294 258458 148350
rect 258278 148170 258334 148226
rect 258402 148170 258458 148226
rect 258278 148046 258334 148102
rect 258402 148046 258458 148102
rect 258278 147922 258334 147978
rect 258402 147922 258458 147978
rect 288998 148294 289054 148350
rect 289122 148294 289178 148350
rect 288998 148170 289054 148226
rect 289122 148170 289178 148226
rect 288998 148046 289054 148102
rect 289122 148046 289178 148102
rect 288998 147922 289054 147978
rect 289122 147922 289178 147978
rect 319718 148294 319774 148350
rect 319842 148294 319898 148350
rect 319718 148170 319774 148226
rect 319842 148170 319898 148226
rect 319718 148046 319774 148102
rect 319842 148046 319898 148102
rect 319718 147922 319774 147978
rect 319842 147922 319898 147978
rect 350438 148294 350494 148350
rect 350562 148294 350618 148350
rect 350438 148170 350494 148226
rect 350562 148170 350618 148226
rect 350438 148046 350494 148102
rect 350562 148046 350618 148102
rect 350438 147922 350494 147978
rect 350562 147922 350618 147978
rect 381158 148294 381214 148350
rect 381282 148294 381338 148350
rect 381158 148170 381214 148226
rect 381282 148170 381338 148226
rect 381158 148046 381214 148102
rect 381282 148046 381338 148102
rect 381158 147922 381214 147978
rect 381282 147922 381338 147978
rect 411878 148294 411934 148350
rect 412002 148294 412058 148350
rect 411878 148170 411934 148226
rect 412002 148170 412058 148226
rect 411878 148046 411934 148102
rect 412002 148046 412058 148102
rect 411878 147922 411934 147978
rect 412002 147922 412058 147978
rect 442598 148294 442654 148350
rect 442722 148294 442778 148350
rect 442598 148170 442654 148226
rect 442722 148170 442778 148226
rect 442598 148046 442654 148102
rect 442722 148046 442778 148102
rect 442598 147922 442654 147978
rect 442722 147922 442778 147978
rect 473318 148294 473374 148350
rect 473442 148294 473498 148350
rect 473318 148170 473374 148226
rect 473442 148170 473498 148226
rect 473318 148046 473374 148102
rect 473442 148046 473498 148102
rect 473318 147922 473374 147978
rect 473442 147922 473498 147978
rect 504038 148294 504094 148350
rect 504162 148294 504218 148350
rect 504038 148170 504094 148226
rect 504162 148170 504218 148226
rect 504038 148046 504094 148102
rect 504162 148046 504218 148102
rect 504038 147922 504094 147978
rect 504162 147922 504218 147978
rect 534758 148294 534814 148350
rect 534882 148294 534938 148350
rect 534758 148170 534814 148226
rect 534882 148170 534938 148226
rect 534758 148046 534814 148102
rect 534882 148046 534938 148102
rect 534758 147922 534814 147978
rect 534882 147922 534938 147978
rect 565478 148294 565534 148350
rect 565602 148294 565658 148350
rect 565478 148170 565534 148226
rect 565602 148170 565658 148226
rect 565478 148046 565534 148102
rect 565602 148046 565658 148102
rect 565478 147922 565534 147978
rect 565602 147922 565658 147978
rect 589194 166294 589250 166350
rect 589318 166294 589374 166350
rect 589442 166294 589498 166350
rect 589566 166294 589622 166350
rect 589194 166170 589250 166226
rect 589318 166170 589374 166226
rect 589442 166170 589498 166226
rect 589566 166170 589622 166226
rect 589194 166046 589250 166102
rect 589318 166046 589374 166102
rect 589442 166046 589498 166102
rect 589566 166046 589622 166102
rect 589194 165922 589250 165978
rect 589318 165922 589374 165978
rect 589442 165922 589498 165978
rect 589566 165922 589622 165978
rect 27878 136294 27934 136350
rect 28002 136294 28058 136350
rect 27878 136170 27934 136226
rect 28002 136170 28058 136226
rect 27878 136046 27934 136102
rect 28002 136046 28058 136102
rect 27878 135922 27934 135978
rect 28002 135922 28058 135978
rect 58598 136294 58654 136350
rect 58722 136294 58778 136350
rect 58598 136170 58654 136226
rect 58722 136170 58778 136226
rect 58598 136046 58654 136102
rect 58722 136046 58778 136102
rect 58598 135922 58654 135978
rect 58722 135922 58778 135978
rect 89318 136294 89374 136350
rect 89442 136294 89498 136350
rect 89318 136170 89374 136226
rect 89442 136170 89498 136226
rect 89318 136046 89374 136102
rect 89442 136046 89498 136102
rect 89318 135922 89374 135978
rect 89442 135922 89498 135978
rect 120038 136294 120094 136350
rect 120162 136294 120218 136350
rect 120038 136170 120094 136226
rect 120162 136170 120218 136226
rect 120038 136046 120094 136102
rect 120162 136046 120218 136102
rect 120038 135922 120094 135978
rect 120162 135922 120218 135978
rect 150758 136294 150814 136350
rect 150882 136294 150938 136350
rect 150758 136170 150814 136226
rect 150882 136170 150938 136226
rect 150758 136046 150814 136102
rect 150882 136046 150938 136102
rect 150758 135922 150814 135978
rect 150882 135922 150938 135978
rect 181478 136294 181534 136350
rect 181602 136294 181658 136350
rect 181478 136170 181534 136226
rect 181602 136170 181658 136226
rect 181478 136046 181534 136102
rect 181602 136046 181658 136102
rect 181478 135922 181534 135978
rect 181602 135922 181658 135978
rect 212198 136294 212254 136350
rect 212322 136294 212378 136350
rect 212198 136170 212254 136226
rect 212322 136170 212378 136226
rect 212198 136046 212254 136102
rect 212322 136046 212378 136102
rect 212198 135922 212254 135978
rect 212322 135922 212378 135978
rect 242918 136294 242974 136350
rect 243042 136294 243098 136350
rect 242918 136170 242974 136226
rect 243042 136170 243098 136226
rect 242918 136046 242974 136102
rect 243042 136046 243098 136102
rect 242918 135922 242974 135978
rect 243042 135922 243098 135978
rect 273638 136294 273694 136350
rect 273762 136294 273818 136350
rect 273638 136170 273694 136226
rect 273762 136170 273818 136226
rect 273638 136046 273694 136102
rect 273762 136046 273818 136102
rect 273638 135922 273694 135978
rect 273762 135922 273818 135978
rect 304358 136294 304414 136350
rect 304482 136294 304538 136350
rect 304358 136170 304414 136226
rect 304482 136170 304538 136226
rect 304358 136046 304414 136102
rect 304482 136046 304538 136102
rect 304358 135922 304414 135978
rect 304482 135922 304538 135978
rect 335078 136294 335134 136350
rect 335202 136294 335258 136350
rect 335078 136170 335134 136226
rect 335202 136170 335258 136226
rect 335078 136046 335134 136102
rect 335202 136046 335258 136102
rect 335078 135922 335134 135978
rect 335202 135922 335258 135978
rect 365798 136294 365854 136350
rect 365922 136294 365978 136350
rect 365798 136170 365854 136226
rect 365922 136170 365978 136226
rect 365798 136046 365854 136102
rect 365922 136046 365978 136102
rect 365798 135922 365854 135978
rect 365922 135922 365978 135978
rect 396518 136294 396574 136350
rect 396642 136294 396698 136350
rect 396518 136170 396574 136226
rect 396642 136170 396698 136226
rect 396518 136046 396574 136102
rect 396642 136046 396698 136102
rect 396518 135922 396574 135978
rect 396642 135922 396698 135978
rect 427238 136294 427294 136350
rect 427362 136294 427418 136350
rect 427238 136170 427294 136226
rect 427362 136170 427418 136226
rect 427238 136046 427294 136102
rect 427362 136046 427418 136102
rect 427238 135922 427294 135978
rect 427362 135922 427418 135978
rect 457958 136294 458014 136350
rect 458082 136294 458138 136350
rect 457958 136170 458014 136226
rect 458082 136170 458138 136226
rect 457958 136046 458014 136102
rect 458082 136046 458138 136102
rect 457958 135922 458014 135978
rect 458082 135922 458138 135978
rect 488678 136294 488734 136350
rect 488802 136294 488858 136350
rect 488678 136170 488734 136226
rect 488802 136170 488858 136226
rect 488678 136046 488734 136102
rect 488802 136046 488858 136102
rect 488678 135922 488734 135978
rect 488802 135922 488858 135978
rect 519398 136294 519454 136350
rect 519522 136294 519578 136350
rect 519398 136170 519454 136226
rect 519522 136170 519578 136226
rect 519398 136046 519454 136102
rect 519522 136046 519578 136102
rect 519398 135922 519454 135978
rect 519522 135922 519578 135978
rect 550118 136294 550174 136350
rect 550242 136294 550298 136350
rect 550118 136170 550174 136226
rect 550242 136170 550298 136226
rect 550118 136046 550174 136102
rect 550242 136046 550298 136102
rect 550118 135922 550174 135978
rect 550242 135922 550298 135978
rect 589194 148294 589250 148350
rect 589318 148294 589374 148350
rect 589442 148294 589498 148350
rect 589566 148294 589622 148350
rect 589194 148170 589250 148226
rect 589318 148170 589374 148226
rect 589442 148170 589498 148226
rect 589566 148170 589622 148226
rect 589194 148046 589250 148102
rect 589318 148046 589374 148102
rect 589442 148046 589498 148102
rect 589566 148046 589622 148102
rect 589194 147922 589250 147978
rect 589318 147922 589374 147978
rect 589442 147922 589498 147978
rect 589566 147922 589622 147978
rect 5514 130294 5570 130350
rect 5638 130294 5694 130350
rect 5762 130294 5818 130350
rect 5886 130294 5942 130350
rect 5514 130170 5570 130226
rect 5638 130170 5694 130226
rect 5762 130170 5818 130226
rect 5886 130170 5942 130226
rect 5514 130046 5570 130102
rect 5638 130046 5694 130102
rect 5762 130046 5818 130102
rect 5886 130046 5942 130102
rect 5514 129922 5570 129978
rect 5638 129922 5694 129978
rect 5762 129922 5818 129978
rect 5886 129922 5942 129978
rect -860 112294 -804 112350
rect -736 112294 -680 112350
rect -612 112294 -556 112350
rect -488 112294 -432 112350
rect -860 112170 -804 112226
rect -736 112170 -680 112226
rect -612 112170 -556 112226
rect -488 112170 -432 112226
rect -860 112046 -804 112102
rect -736 112046 -680 112102
rect -612 112046 -556 112102
rect -488 112046 -432 112102
rect -860 111922 -804 111978
rect -736 111922 -680 111978
rect -612 111922 -556 111978
rect -488 111922 -432 111978
rect 12518 130294 12574 130350
rect 12642 130294 12698 130350
rect 12518 130170 12574 130226
rect 12642 130170 12698 130226
rect 12518 130046 12574 130102
rect 12642 130046 12698 130102
rect 12518 129922 12574 129978
rect 12642 129922 12698 129978
rect 43238 130294 43294 130350
rect 43362 130294 43418 130350
rect 43238 130170 43294 130226
rect 43362 130170 43418 130226
rect 43238 130046 43294 130102
rect 43362 130046 43418 130102
rect 43238 129922 43294 129978
rect 43362 129922 43418 129978
rect 73958 130294 74014 130350
rect 74082 130294 74138 130350
rect 73958 130170 74014 130226
rect 74082 130170 74138 130226
rect 73958 130046 74014 130102
rect 74082 130046 74138 130102
rect 73958 129922 74014 129978
rect 74082 129922 74138 129978
rect 104678 130294 104734 130350
rect 104802 130294 104858 130350
rect 104678 130170 104734 130226
rect 104802 130170 104858 130226
rect 104678 130046 104734 130102
rect 104802 130046 104858 130102
rect 104678 129922 104734 129978
rect 104802 129922 104858 129978
rect 135398 130294 135454 130350
rect 135522 130294 135578 130350
rect 135398 130170 135454 130226
rect 135522 130170 135578 130226
rect 135398 130046 135454 130102
rect 135522 130046 135578 130102
rect 135398 129922 135454 129978
rect 135522 129922 135578 129978
rect 166118 130294 166174 130350
rect 166242 130294 166298 130350
rect 166118 130170 166174 130226
rect 166242 130170 166298 130226
rect 166118 130046 166174 130102
rect 166242 130046 166298 130102
rect 166118 129922 166174 129978
rect 166242 129922 166298 129978
rect 196838 130294 196894 130350
rect 196962 130294 197018 130350
rect 196838 130170 196894 130226
rect 196962 130170 197018 130226
rect 196838 130046 196894 130102
rect 196962 130046 197018 130102
rect 196838 129922 196894 129978
rect 196962 129922 197018 129978
rect 227558 130294 227614 130350
rect 227682 130294 227738 130350
rect 227558 130170 227614 130226
rect 227682 130170 227738 130226
rect 227558 130046 227614 130102
rect 227682 130046 227738 130102
rect 227558 129922 227614 129978
rect 227682 129922 227738 129978
rect 258278 130294 258334 130350
rect 258402 130294 258458 130350
rect 258278 130170 258334 130226
rect 258402 130170 258458 130226
rect 258278 130046 258334 130102
rect 258402 130046 258458 130102
rect 258278 129922 258334 129978
rect 258402 129922 258458 129978
rect 288998 130294 289054 130350
rect 289122 130294 289178 130350
rect 288998 130170 289054 130226
rect 289122 130170 289178 130226
rect 288998 130046 289054 130102
rect 289122 130046 289178 130102
rect 288998 129922 289054 129978
rect 289122 129922 289178 129978
rect 319718 130294 319774 130350
rect 319842 130294 319898 130350
rect 319718 130170 319774 130226
rect 319842 130170 319898 130226
rect 319718 130046 319774 130102
rect 319842 130046 319898 130102
rect 319718 129922 319774 129978
rect 319842 129922 319898 129978
rect 350438 130294 350494 130350
rect 350562 130294 350618 130350
rect 350438 130170 350494 130226
rect 350562 130170 350618 130226
rect 350438 130046 350494 130102
rect 350562 130046 350618 130102
rect 350438 129922 350494 129978
rect 350562 129922 350618 129978
rect 381158 130294 381214 130350
rect 381282 130294 381338 130350
rect 381158 130170 381214 130226
rect 381282 130170 381338 130226
rect 381158 130046 381214 130102
rect 381282 130046 381338 130102
rect 381158 129922 381214 129978
rect 381282 129922 381338 129978
rect 411878 130294 411934 130350
rect 412002 130294 412058 130350
rect 411878 130170 411934 130226
rect 412002 130170 412058 130226
rect 411878 130046 411934 130102
rect 412002 130046 412058 130102
rect 411878 129922 411934 129978
rect 412002 129922 412058 129978
rect 442598 130294 442654 130350
rect 442722 130294 442778 130350
rect 442598 130170 442654 130226
rect 442722 130170 442778 130226
rect 442598 130046 442654 130102
rect 442722 130046 442778 130102
rect 442598 129922 442654 129978
rect 442722 129922 442778 129978
rect 473318 130294 473374 130350
rect 473442 130294 473498 130350
rect 473318 130170 473374 130226
rect 473442 130170 473498 130226
rect 473318 130046 473374 130102
rect 473442 130046 473498 130102
rect 473318 129922 473374 129978
rect 473442 129922 473498 129978
rect 504038 130294 504094 130350
rect 504162 130294 504218 130350
rect 504038 130170 504094 130226
rect 504162 130170 504218 130226
rect 504038 130046 504094 130102
rect 504162 130046 504218 130102
rect 504038 129922 504094 129978
rect 504162 129922 504218 129978
rect 534758 130294 534814 130350
rect 534882 130294 534938 130350
rect 534758 130170 534814 130226
rect 534882 130170 534938 130226
rect 534758 130046 534814 130102
rect 534882 130046 534938 130102
rect 534758 129922 534814 129978
rect 534882 129922 534938 129978
rect 565478 130294 565534 130350
rect 565602 130294 565658 130350
rect 565478 130170 565534 130226
rect 565602 130170 565658 130226
rect 565478 130046 565534 130102
rect 565602 130046 565658 130102
rect 565478 129922 565534 129978
rect 565602 129922 565658 129978
rect 592914 208294 592970 208350
rect 593038 208294 593094 208350
rect 593162 208294 593218 208350
rect 593286 208294 593342 208350
rect 592914 208170 592970 208226
rect 593038 208170 593094 208226
rect 593162 208170 593218 208226
rect 593286 208170 593342 208226
rect 592914 208046 592970 208102
rect 593038 208046 593094 208102
rect 593162 208046 593218 208102
rect 593286 208046 593342 208102
rect 592914 207922 592970 207978
rect 593038 207922 593094 207978
rect 593162 207922 593218 207978
rect 593286 207922 593342 207978
rect 592914 190294 592970 190350
rect 593038 190294 593094 190350
rect 593162 190294 593218 190350
rect 593286 190294 593342 190350
rect 592914 190170 592970 190226
rect 593038 190170 593094 190226
rect 593162 190170 593218 190226
rect 593286 190170 593342 190226
rect 592914 190046 592970 190102
rect 593038 190046 593094 190102
rect 593162 190046 593218 190102
rect 593286 190046 593342 190102
rect 592914 189922 592970 189978
rect 593038 189922 593094 189978
rect 593162 189922 593218 189978
rect 593286 189922 593342 189978
rect 592914 172294 592970 172350
rect 593038 172294 593094 172350
rect 593162 172294 593218 172350
rect 593286 172294 593342 172350
rect 592914 172170 592970 172226
rect 593038 172170 593094 172226
rect 593162 172170 593218 172226
rect 593286 172170 593342 172226
rect 592914 172046 592970 172102
rect 593038 172046 593094 172102
rect 593162 172046 593218 172102
rect 593286 172046 593342 172102
rect 592914 171922 592970 171978
rect 593038 171922 593094 171978
rect 593162 171922 593218 171978
rect 593286 171922 593342 171978
rect 592914 154294 592970 154350
rect 593038 154294 593094 154350
rect 593162 154294 593218 154350
rect 593286 154294 593342 154350
rect 592914 154170 592970 154226
rect 593038 154170 593094 154226
rect 593162 154170 593218 154226
rect 593286 154170 593342 154226
rect 592914 154046 592970 154102
rect 593038 154046 593094 154102
rect 593162 154046 593218 154102
rect 593286 154046 593342 154102
rect 592914 153922 592970 153978
rect 593038 153922 593094 153978
rect 593162 153922 593218 153978
rect 593286 153922 593342 153978
rect 589194 130294 589250 130350
rect 589318 130294 589374 130350
rect 589442 130294 589498 130350
rect 589566 130294 589622 130350
rect 589194 130170 589250 130226
rect 589318 130170 589374 130226
rect 589442 130170 589498 130226
rect 589566 130170 589622 130226
rect 589194 130046 589250 130102
rect 589318 130046 589374 130102
rect 589442 130046 589498 130102
rect 589566 130046 589622 130102
rect 589194 129922 589250 129978
rect 589318 129922 589374 129978
rect 589442 129922 589498 129978
rect 589566 129922 589622 129978
rect 27878 118294 27934 118350
rect 28002 118294 28058 118350
rect 27878 118170 27934 118226
rect 28002 118170 28058 118226
rect 27878 118046 27934 118102
rect 28002 118046 28058 118102
rect 27878 117922 27934 117978
rect 28002 117922 28058 117978
rect 58598 118294 58654 118350
rect 58722 118294 58778 118350
rect 58598 118170 58654 118226
rect 58722 118170 58778 118226
rect 58598 118046 58654 118102
rect 58722 118046 58778 118102
rect 58598 117922 58654 117978
rect 58722 117922 58778 117978
rect 89318 118294 89374 118350
rect 89442 118294 89498 118350
rect 89318 118170 89374 118226
rect 89442 118170 89498 118226
rect 89318 118046 89374 118102
rect 89442 118046 89498 118102
rect 89318 117922 89374 117978
rect 89442 117922 89498 117978
rect 120038 118294 120094 118350
rect 120162 118294 120218 118350
rect 120038 118170 120094 118226
rect 120162 118170 120218 118226
rect 120038 118046 120094 118102
rect 120162 118046 120218 118102
rect 120038 117922 120094 117978
rect 120162 117922 120218 117978
rect 150758 118294 150814 118350
rect 150882 118294 150938 118350
rect 150758 118170 150814 118226
rect 150882 118170 150938 118226
rect 150758 118046 150814 118102
rect 150882 118046 150938 118102
rect 150758 117922 150814 117978
rect 150882 117922 150938 117978
rect 181478 118294 181534 118350
rect 181602 118294 181658 118350
rect 181478 118170 181534 118226
rect 181602 118170 181658 118226
rect 181478 118046 181534 118102
rect 181602 118046 181658 118102
rect 181478 117922 181534 117978
rect 181602 117922 181658 117978
rect 212198 118294 212254 118350
rect 212322 118294 212378 118350
rect 212198 118170 212254 118226
rect 212322 118170 212378 118226
rect 212198 118046 212254 118102
rect 212322 118046 212378 118102
rect 212198 117922 212254 117978
rect 212322 117922 212378 117978
rect 242918 118294 242974 118350
rect 243042 118294 243098 118350
rect 242918 118170 242974 118226
rect 243042 118170 243098 118226
rect 242918 118046 242974 118102
rect 243042 118046 243098 118102
rect 242918 117922 242974 117978
rect 243042 117922 243098 117978
rect 273638 118294 273694 118350
rect 273762 118294 273818 118350
rect 273638 118170 273694 118226
rect 273762 118170 273818 118226
rect 273638 118046 273694 118102
rect 273762 118046 273818 118102
rect 273638 117922 273694 117978
rect 273762 117922 273818 117978
rect 304358 118294 304414 118350
rect 304482 118294 304538 118350
rect 304358 118170 304414 118226
rect 304482 118170 304538 118226
rect 304358 118046 304414 118102
rect 304482 118046 304538 118102
rect 304358 117922 304414 117978
rect 304482 117922 304538 117978
rect 335078 118294 335134 118350
rect 335202 118294 335258 118350
rect 335078 118170 335134 118226
rect 335202 118170 335258 118226
rect 335078 118046 335134 118102
rect 335202 118046 335258 118102
rect 335078 117922 335134 117978
rect 335202 117922 335258 117978
rect 365798 118294 365854 118350
rect 365922 118294 365978 118350
rect 365798 118170 365854 118226
rect 365922 118170 365978 118226
rect 365798 118046 365854 118102
rect 365922 118046 365978 118102
rect 365798 117922 365854 117978
rect 365922 117922 365978 117978
rect 396518 118294 396574 118350
rect 396642 118294 396698 118350
rect 396518 118170 396574 118226
rect 396642 118170 396698 118226
rect 396518 118046 396574 118102
rect 396642 118046 396698 118102
rect 396518 117922 396574 117978
rect 396642 117922 396698 117978
rect 427238 118294 427294 118350
rect 427362 118294 427418 118350
rect 427238 118170 427294 118226
rect 427362 118170 427418 118226
rect 427238 118046 427294 118102
rect 427362 118046 427418 118102
rect 427238 117922 427294 117978
rect 427362 117922 427418 117978
rect 457958 118294 458014 118350
rect 458082 118294 458138 118350
rect 457958 118170 458014 118226
rect 458082 118170 458138 118226
rect 457958 118046 458014 118102
rect 458082 118046 458138 118102
rect 457958 117922 458014 117978
rect 458082 117922 458138 117978
rect 488678 118294 488734 118350
rect 488802 118294 488858 118350
rect 488678 118170 488734 118226
rect 488802 118170 488858 118226
rect 488678 118046 488734 118102
rect 488802 118046 488858 118102
rect 488678 117922 488734 117978
rect 488802 117922 488858 117978
rect 519398 118294 519454 118350
rect 519522 118294 519578 118350
rect 519398 118170 519454 118226
rect 519522 118170 519578 118226
rect 519398 118046 519454 118102
rect 519522 118046 519578 118102
rect 519398 117922 519454 117978
rect 519522 117922 519578 117978
rect 550118 118294 550174 118350
rect 550242 118294 550298 118350
rect 550118 118170 550174 118226
rect 550242 118170 550298 118226
rect 550118 118046 550174 118102
rect 550242 118046 550298 118102
rect 550118 117922 550174 117978
rect 550242 117922 550298 117978
rect 5514 112294 5570 112350
rect 5638 112294 5694 112350
rect 5762 112294 5818 112350
rect 5886 112294 5942 112350
rect 5514 112170 5570 112226
rect 5638 112170 5694 112226
rect 5762 112170 5818 112226
rect 5886 112170 5942 112226
rect 5514 112046 5570 112102
rect 5638 112046 5694 112102
rect 5762 112046 5818 112102
rect 5886 112046 5942 112102
rect 5514 111922 5570 111978
rect 5638 111922 5694 111978
rect 5762 111922 5818 111978
rect 5886 111922 5942 111978
rect -860 94294 -804 94350
rect -736 94294 -680 94350
rect -612 94294 -556 94350
rect -488 94294 -432 94350
rect -860 94170 -804 94226
rect -736 94170 -680 94226
rect -612 94170 -556 94226
rect -488 94170 -432 94226
rect -860 94046 -804 94102
rect -736 94046 -680 94102
rect -612 94046 -556 94102
rect -488 94046 -432 94102
rect -860 93922 -804 93978
rect -736 93922 -680 93978
rect -612 93922 -556 93978
rect -488 93922 -432 93978
rect 12518 112294 12574 112350
rect 12642 112294 12698 112350
rect 12518 112170 12574 112226
rect 12642 112170 12698 112226
rect 12518 112046 12574 112102
rect 12642 112046 12698 112102
rect 12518 111922 12574 111978
rect 12642 111922 12698 111978
rect 43238 112294 43294 112350
rect 43362 112294 43418 112350
rect 43238 112170 43294 112226
rect 43362 112170 43418 112226
rect 43238 112046 43294 112102
rect 43362 112046 43418 112102
rect 43238 111922 43294 111978
rect 43362 111922 43418 111978
rect 73958 112294 74014 112350
rect 74082 112294 74138 112350
rect 73958 112170 74014 112226
rect 74082 112170 74138 112226
rect 73958 112046 74014 112102
rect 74082 112046 74138 112102
rect 73958 111922 74014 111978
rect 74082 111922 74138 111978
rect 104678 112294 104734 112350
rect 104802 112294 104858 112350
rect 104678 112170 104734 112226
rect 104802 112170 104858 112226
rect 104678 112046 104734 112102
rect 104802 112046 104858 112102
rect 104678 111922 104734 111978
rect 104802 111922 104858 111978
rect 135398 112294 135454 112350
rect 135522 112294 135578 112350
rect 135398 112170 135454 112226
rect 135522 112170 135578 112226
rect 135398 112046 135454 112102
rect 135522 112046 135578 112102
rect 135398 111922 135454 111978
rect 135522 111922 135578 111978
rect 166118 112294 166174 112350
rect 166242 112294 166298 112350
rect 166118 112170 166174 112226
rect 166242 112170 166298 112226
rect 166118 112046 166174 112102
rect 166242 112046 166298 112102
rect 166118 111922 166174 111978
rect 166242 111922 166298 111978
rect 196838 112294 196894 112350
rect 196962 112294 197018 112350
rect 196838 112170 196894 112226
rect 196962 112170 197018 112226
rect 196838 112046 196894 112102
rect 196962 112046 197018 112102
rect 196838 111922 196894 111978
rect 196962 111922 197018 111978
rect 227558 112294 227614 112350
rect 227682 112294 227738 112350
rect 227558 112170 227614 112226
rect 227682 112170 227738 112226
rect 227558 112046 227614 112102
rect 227682 112046 227738 112102
rect 227558 111922 227614 111978
rect 227682 111922 227738 111978
rect 258278 112294 258334 112350
rect 258402 112294 258458 112350
rect 258278 112170 258334 112226
rect 258402 112170 258458 112226
rect 258278 112046 258334 112102
rect 258402 112046 258458 112102
rect 258278 111922 258334 111978
rect 258402 111922 258458 111978
rect 288998 112294 289054 112350
rect 289122 112294 289178 112350
rect 288998 112170 289054 112226
rect 289122 112170 289178 112226
rect 288998 112046 289054 112102
rect 289122 112046 289178 112102
rect 288998 111922 289054 111978
rect 289122 111922 289178 111978
rect 319718 112294 319774 112350
rect 319842 112294 319898 112350
rect 319718 112170 319774 112226
rect 319842 112170 319898 112226
rect 319718 112046 319774 112102
rect 319842 112046 319898 112102
rect 319718 111922 319774 111978
rect 319842 111922 319898 111978
rect 350438 112294 350494 112350
rect 350562 112294 350618 112350
rect 350438 112170 350494 112226
rect 350562 112170 350618 112226
rect 350438 112046 350494 112102
rect 350562 112046 350618 112102
rect 350438 111922 350494 111978
rect 350562 111922 350618 111978
rect 381158 112294 381214 112350
rect 381282 112294 381338 112350
rect 381158 112170 381214 112226
rect 381282 112170 381338 112226
rect 381158 112046 381214 112102
rect 381282 112046 381338 112102
rect 381158 111922 381214 111978
rect 381282 111922 381338 111978
rect 411878 112294 411934 112350
rect 412002 112294 412058 112350
rect 411878 112170 411934 112226
rect 412002 112170 412058 112226
rect 411878 112046 411934 112102
rect 412002 112046 412058 112102
rect 411878 111922 411934 111978
rect 412002 111922 412058 111978
rect 442598 112294 442654 112350
rect 442722 112294 442778 112350
rect 442598 112170 442654 112226
rect 442722 112170 442778 112226
rect 442598 112046 442654 112102
rect 442722 112046 442778 112102
rect 442598 111922 442654 111978
rect 442722 111922 442778 111978
rect 473318 112294 473374 112350
rect 473442 112294 473498 112350
rect 473318 112170 473374 112226
rect 473442 112170 473498 112226
rect 473318 112046 473374 112102
rect 473442 112046 473498 112102
rect 473318 111922 473374 111978
rect 473442 111922 473498 111978
rect 504038 112294 504094 112350
rect 504162 112294 504218 112350
rect 504038 112170 504094 112226
rect 504162 112170 504218 112226
rect 504038 112046 504094 112102
rect 504162 112046 504218 112102
rect 504038 111922 504094 111978
rect 504162 111922 504218 111978
rect 534758 112294 534814 112350
rect 534882 112294 534938 112350
rect 534758 112170 534814 112226
rect 534882 112170 534938 112226
rect 534758 112046 534814 112102
rect 534882 112046 534938 112102
rect 534758 111922 534814 111978
rect 534882 111922 534938 111978
rect 565478 112294 565534 112350
rect 565602 112294 565658 112350
rect 565478 112170 565534 112226
rect 565602 112170 565658 112226
rect 565478 112046 565534 112102
rect 565602 112046 565658 112102
rect 565478 111922 565534 111978
rect 565602 111922 565658 111978
rect 592914 136294 592970 136350
rect 593038 136294 593094 136350
rect 593162 136294 593218 136350
rect 593286 136294 593342 136350
rect 592914 136170 592970 136226
rect 593038 136170 593094 136226
rect 593162 136170 593218 136226
rect 593286 136170 593342 136226
rect 592914 136046 592970 136102
rect 593038 136046 593094 136102
rect 593162 136046 593218 136102
rect 593286 136046 593342 136102
rect 592914 135922 592970 135978
rect 593038 135922 593094 135978
rect 593162 135922 593218 135978
rect 593286 135922 593342 135978
rect 592914 118294 592970 118350
rect 593038 118294 593094 118350
rect 593162 118294 593218 118350
rect 593286 118294 593342 118350
rect 592914 118170 592970 118226
rect 593038 118170 593094 118226
rect 593162 118170 593218 118226
rect 593286 118170 593342 118226
rect 592914 118046 592970 118102
rect 593038 118046 593094 118102
rect 593162 118046 593218 118102
rect 593286 118046 593342 118102
rect 592914 117922 592970 117978
rect 593038 117922 593094 117978
rect 593162 117922 593218 117978
rect 593286 117922 593342 117978
rect 589194 112294 589250 112350
rect 589318 112294 589374 112350
rect 589442 112294 589498 112350
rect 589566 112294 589622 112350
rect 589194 112170 589250 112226
rect 589318 112170 589374 112226
rect 589442 112170 589498 112226
rect 589566 112170 589622 112226
rect 589194 112046 589250 112102
rect 589318 112046 589374 112102
rect 589442 112046 589498 112102
rect 589566 112046 589622 112102
rect 589194 111922 589250 111978
rect 589318 111922 589374 111978
rect 589442 111922 589498 111978
rect 589566 111922 589622 111978
rect 5514 94294 5570 94350
rect 5638 94294 5694 94350
rect 5762 94294 5818 94350
rect 5886 94294 5942 94350
rect 5514 94170 5570 94226
rect 5638 94170 5694 94226
rect 5762 94170 5818 94226
rect 5886 94170 5942 94226
rect 5514 94046 5570 94102
rect 5638 94046 5694 94102
rect 5762 94046 5818 94102
rect 5886 94046 5942 94102
rect 5514 93922 5570 93978
rect 5638 93922 5694 93978
rect 5762 93922 5818 93978
rect 5886 93922 5942 93978
rect -860 76294 -804 76350
rect -736 76294 -680 76350
rect -612 76294 -556 76350
rect -488 76294 -432 76350
rect -860 76170 -804 76226
rect -736 76170 -680 76226
rect -612 76170 -556 76226
rect -488 76170 -432 76226
rect -860 76046 -804 76102
rect -736 76046 -680 76102
rect -612 76046 -556 76102
rect -488 76046 -432 76102
rect -860 75922 -804 75978
rect -736 75922 -680 75978
rect -612 75922 -556 75978
rect -488 75922 -432 75978
rect 27878 100294 27934 100350
rect 28002 100294 28058 100350
rect 27878 100170 27934 100226
rect 28002 100170 28058 100226
rect 27878 100046 27934 100102
rect 28002 100046 28058 100102
rect 27878 99922 27934 99978
rect 28002 99922 28058 99978
rect 58598 100294 58654 100350
rect 58722 100294 58778 100350
rect 58598 100170 58654 100226
rect 58722 100170 58778 100226
rect 58598 100046 58654 100102
rect 58722 100046 58778 100102
rect 58598 99922 58654 99978
rect 58722 99922 58778 99978
rect 89318 100294 89374 100350
rect 89442 100294 89498 100350
rect 89318 100170 89374 100226
rect 89442 100170 89498 100226
rect 89318 100046 89374 100102
rect 89442 100046 89498 100102
rect 89318 99922 89374 99978
rect 89442 99922 89498 99978
rect 120038 100294 120094 100350
rect 120162 100294 120218 100350
rect 120038 100170 120094 100226
rect 120162 100170 120218 100226
rect 120038 100046 120094 100102
rect 120162 100046 120218 100102
rect 120038 99922 120094 99978
rect 120162 99922 120218 99978
rect 150758 100294 150814 100350
rect 150882 100294 150938 100350
rect 150758 100170 150814 100226
rect 150882 100170 150938 100226
rect 150758 100046 150814 100102
rect 150882 100046 150938 100102
rect 150758 99922 150814 99978
rect 150882 99922 150938 99978
rect 181478 100294 181534 100350
rect 181602 100294 181658 100350
rect 181478 100170 181534 100226
rect 181602 100170 181658 100226
rect 181478 100046 181534 100102
rect 181602 100046 181658 100102
rect 181478 99922 181534 99978
rect 181602 99922 181658 99978
rect 212198 100294 212254 100350
rect 212322 100294 212378 100350
rect 212198 100170 212254 100226
rect 212322 100170 212378 100226
rect 212198 100046 212254 100102
rect 212322 100046 212378 100102
rect 212198 99922 212254 99978
rect 212322 99922 212378 99978
rect 242918 100294 242974 100350
rect 243042 100294 243098 100350
rect 242918 100170 242974 100226
rect 243042 100170 243098 100226
rect 242918 100046 242974 100102
rect 243042 100046 243098 100102
rect 242918 99922 242974 99978
rect 243042 99922 243098 99978
rect 273638 100294 273694 100350
rect 273762 100294 273818 100350
rect 273638 100170 273694 100226
rect 273762 100170 273818 100226
rect 273638 100046 273694 100102
rect 273762 100046 273818 100102
rect 273638 99922 273694 99978
rect 273762 99922 273818 99978
rect 304358 100294 304414 100350
rect 304482 100294 304538 100350
rect 304358 100170 304414 100226
rect 304482 100170 304538 100226
rect 304358 100046 304414 100102
rect 304482 100046 304538 100102
rect 304358 99922 304414 99978
rect 304482 99922 304538 99978
rect 335078 100294 335134 100350
rect 335202 100294 335258 100350
rect 335078 100170 335134 100226
rect 335202 100170 335258 100226
rect 335078 100046 335134 100102
rect 335202 100046 335258 100102
rect 335078 99922 335134 99978
rect 335202 99922 335258 99978
rect 365798 100294 365854 100350
rect 365922 100294 365978 100350
rect 365798 100170 365854 100226
rect 365922 100170 365978 100226
rect 365798 100046 365854 100102
rect 365922 100046 365978 100102
rect 365798 99922 365854 99978
rect 365922 99922 365978 99978
rect 396518 100294 396574 100350
rect 396642 100294 396698 100350
rect 396518 100170 396574 100226
rect 396642 100170 396698 100226
rect 396518 100046 396574 100102
rect 396642 100046 396698 100102
rect 396518 99922 396574 99978
rect 396642 99922 396698 99978
rect 427238 100294 427294 100350
rect 427362 100294 427418 100350
rect 427238 100170 427294 100226
rect 427362 100170 427418 100226
rect 427238 100046 427294 100102
rect 427362 100046 427418 100102
rect 427238 99922 427294 99978
rect 427362 99922 427418 99978
rect 457958 100294 458014 100350
rect 458082 100294 458138 100350
rect 457958 100170 458014 100226
rect 458082 100170 458138 100226
rect 457958 100046 458014 100102
rect 458082 100046 458138 100102
rect 457958 99922 458014 99978
rect 458082 99922 458138 99978
rect 488678 100294 488734 100350
rect 488802 100294 488858 100350
rect 488678 100170 488734 100226
rect 488802 100170 488858 100226
rect 488678 100046 488734 100102
rect 488802 100046 488858 100102
rect 488678 99922 488734 99978
rect 488802 99922 488858 99978
rect 519398 100294 519454 100350
rect 519522 100294 519578 100350
rect 519398 100170 519454 100226
rect 519522 100170 519578 100226
rect 519398 100046 519454 100102
rect 519522 100046 519578 100102
rect 519398 99922 519454 99978
rect 519522 99922 519578 99978
rect 550118 100294 550174 100350
rect 550242 100294 550298 100350
rect 550118 100170 550174 100226
rect 550242 100170 550298 100226
rect 550118 100046 550174 100102
rect 550242 100046 550298 100102
rect 550118 99922 550174 99978
rect 550242 99922 550298 99978
rect 12518 94294 12574 94350
rect 12642 94294 12698 94350
rect 12518 94170 12574 94226
rect 12642 94170 12698 94226
rect 12518 94046 12574 94102
rect 12642 94046 12698 94102
rect 12518 93922 12574 93978
rect 12642 93922 12698 93978
rect 43238 94294 43294 94350
rect 43362 94294 43418 94350
rect 43238 94170 43294 94226
rect 43362 94170 43418 94226
rect 43238 94046 43294 94102
rect 43362 94046 43418 94102
rect 43238 93922 43294 93978
rect 43362 93922 43418 93978
rect 73958 94294 74014 94350
rect 74082 94294 74138 94350
rect 73958 94170 74014 94226
rect 74082 94170 74138 94226
rect 73958 94046 74014 94102
rect 74082 94046 74138 94102
rect 73958 93922 74014 93978
rect 74082 93922 74138 93978
rect 104678 94294 104734 94350
rect 104802 94294 104858 94350
rect 104678 94170 104734 94226
rect 104802 94170 104858 94226
rect 104678 94046 104734 94102
rect 104802 94046 104858 94102
rect 104678 93922 104734 93978
rect 104802 93922 104858 93978
rect 135398 94294 135454 94350
rect 135522 94294 135578 94350
rect 135398 94170 135454 94226
rect 135522 94170 135578 94226
rect 135398 94046 135454 94102
rect 135522 94046 135578 94102
rect 135398 93922 135454 93978
rect 135522 93922 135578 93978
rect 166118 94294 166174 94350
rect 166242 94294 166298 94350
rect 166118 94170 166174 94226
rect 166242 94170 166298 94226
rect 166118 94046 166174 94102
rect 166242 94046 166298 94102
rect 166118 93922 166174 93978
rect 166242 93922 166298 93978
rect 196838 94294 196894 94350
rect 196962 94294 197018 94350
rect 196838 94170 196894 94226
rect 196962 94170 197018 94226
rect 196838 94046 196894 94102
rect 196962 94046 197018 94102
rect 196838 93922 196894 93978
rect 196962 93922 197018 93978
rect 227558 94294 227614 94350
rect 227682 94294 227738 94350
rect 227558 94170 227614 94226
rect 227682 94170 227738 94226
rect 227558 94046 227614 94102
rect 227682 94046 227738 94102
rect 227558 93922 227614 93978
rect 227682 93922 227738 93978
rect 258278 94294 258334 94350
rect 258402 94294 258458 94350
rect 258278 94170 258334 94226
rect 258402 94170 258458 94226
rect 258278 94046 258334 94102
rect 258402 94046 258458 94102
rect 258278 93922 258334 93978
rect 258402 93922 258458 93978
rect 288998 94294 289054 94350
rect 289122 94294 289178 94350
rect 288998 94170 289054 94226
rect 289122 94170 289178 94226
rect 288998 94046 289054 94102
rect 289122 94046 289178 94102
rect 288998 93922 289054 93978
rect 289122 93922 289178 93978
rect 319718 94294 319774 94350
rect 319842 94294 319898 94350
rect 319718 94170 319774 94226
rect 319842 94170 319898 94226
rect 319718 94046 319774 94102
rect 319842 94046 319898 94102
rect 319718 93922 319774 93978
rect 319842 93922 319898 93978
rect 350438 94294 350494 94350
rect 350562 94294 350618 94350
rect 350438 94170 350494 94226
rect 350562 94170 350618 94226
rect 350438 94046 350494 94102
rect 350562 94046 350618 94102
rect 350438 93922 350494 93978
rect 350562 93922 350618 93978
rect 381158 94294 381214 94350
rect 381282 94294 381338 94350
rect 381158 94170 381214 94226
rect 381282 94170 381338 94226
rect 381158 94046 381214 94102
rect 381282 94046 381338 94102
rect 381158 93922 381214 93978
rect 381282 93922 381338 93978
rect 411878 94294 411934 94350
rect 412002 94294 412058 94350
rect 411878 94170 411934 94226
rect 412002 94170 412058 94226
rect 411878 94046 411934 94102
rect 412002 94046 412058 94102
rect 411878 93922 411934 93978
rect 412002 93922 412058 93978
rect 442598 94294 442654 94350
rect 442722 94294 442778 94350
rect 442598 94170 442654 94226
rect 442722 94170 442778 94226
rect 442598 94046 442654 94102
rect 442722 94046 442778 94102
rect 442598 93922 442654 93978
rect 442722 93922 442778 93978
rect 473318 94294 473374 94350
rect 473442 94294 473498 94350
rect 473318 94170 473374 94226
rect 473442 94170 473498 94226
rect 473318 94046 473374 94102
rect 473442 94046 473498 94102
rect 473318 93922 473374 93978
rect 473442 93922 473498 93978
rect 504038 94294 504094 94350
rect 504162 94294 504218 94350
rect 504038 94170 504094 94226
rect 504162 94170 504218 94226
rect 504038 94046 504094 94102
rect 504162 94046 504218 94102
rect 504038 93922 504094 93978
rect 504162 93922 504218 93978
rect 534758 94294 534814 94350
rect 534882 94294 534938 94350
rect 534758 94170 534814 94226
rect 534882 94170 534938 94226
rect 534758 94046 534814 94102
rect 534882 94046 534938 94102
rect 534758 93922 534814 93978
rect 534882 93922 534938 93978
rect 565478 94294 565534 94350
rect 565602 94294 565658 94350
rect 565478 94170 565534 94226
rect 565602 94170 565658 94226
rect 565478 94046 565534 94102
rect 565602 94046 565658 94102
rect 565478 93922 565534 93978
rect 565602 93922 565658 93978
rect 589194 94294 589250 94350
rect 589318 94294 589374 94350
rect 589442 94294 589498 94350
rect 589566 94294 589622 94350
rect 589194 94170 589250 94226
rect 589318 94170 589374 94226
rect 589442 94170 589498 94226
rect 589566 94170 589622 94226
rect 589194 94046 589250 94102
rect 589318 94046 589374 94102
rect 589442 94046 589498 94102
rect 589566 94046 589622 94102
rect 589194 93922 589250 93978
rect 589318 93922 589374 93978
rect 589442 93922 589498 93978
rect 589566 93922 589622 93978
rect 27878 82294 27934 82350
rect 28002 82294 28058 82350
rect 27878 82170 27934 82226
rect 28002 82170 28058 82226
rect 27878 82046 27934 82102
rect 28002 82046 28058 82102
rect 27878 81922 27934 81978
rect 28002 81922 28058 81978
rect 58598 82294 58654 82350
rect 58722 82294 58778 82350
rect 58598 82170 58654 82226
rect 58722 82170 58778 82226
rect 58598 82046 58654 82102
rect 58722 82046 58778 82102
rect 58598 81922 58654 81978
rect 58722 81922 58778 81978
rect 89318 82294 89374 82350
rect 89442 82294 89498 82350
rect 89318 82170 89374 82226
rect 89442 82170 89498 82226
rect 89318 82046 89374 82102
rect 89442 82046 89498 82102
rect 89318 81922 89374 81978
rect 89442 81922 89498 81978
rect 120038 82294 120094 82350
rect 120162 82294 120218 82350
rect 120038 82170 120094 82226
rect 120162 82170 120218 82226
rect 120038 82046 120094 82102
rect 120162 82046 120218 82102
rect 120038 81922 120094 81978
rect 120162 81922 120218 81978
rect 150758 82294 150814 82350
rect 150882 82294 150938 82350
rect 150758 82170 150814 82226
rect 150882 82170 150938 82226
rect 150758 82046 150814 82102
rect 150882 82046 150938 82102
rect 150758 81922 150814 81978
rect 150882 81922 150938 81978
rect 181478 82294 181534 82350
rect 181602 82294 181658 82350
rect 181478 82170 181534 82226
rect 181602 82170 181658 82226
rect 181478 82046 181534 82102
rect 181602 82046 181658 82102
rect 181478 81922 181534 81978
rect 181602 81922 181658 81978
rect 212198 82294 212254 82350
rect 212322 82294 212378 82350
rect 212198 82170 212254 82226
rect 212322 82170 212378 82226
rect 212198 82046 212254 82102
rect 212322 82046 212378 82102
rect 212198 81922 212254 81978
rect 212322 81922 212378 81978
rect 242918 82294 242974 82350
rect 243042 82294 243098 82350
rect 242918 82170 242974 82226
rect 243042 82170 243098 82226
rect 242918 82046 242974 82102
rect 243042 82046 243098 82102
rect 242918 81922 242974 81978
rect 243042 81922 243098 81978
rect 273638 82294 273694 82350
rect 273762 82294 273818 82350
rect 273638 82170 273694 82226
rect 273762 82170 273818 82226
rect 273638 82046 273694 82102
rect 273762 82046 273818 82102
rect 273638 81922 273694 81978
rect 273762 81922 273818 81978
rect 304358 82294 304414 82350
rect 304482 82294 304538 82350
rect 304358 82170 304414 82226
rect 304482 82170 304538 82226
rect 304358 82046 304414 82102
rect 304482 82046 304538 82102
rect 304358 81922 304414 81978
rect 304482 81922 304538 81978
rect 335078 82294 335134 82350
rect 335202 82294 335258 82350
rect 335078 82170 335134 82226
rect 335202 82170 335258 82226
rect 335078 82046 335134 82102
rect 335202 82046 335258 82102
rect 335078 81922 335134 81978
rect 335202 81922 335258 81978
rect 365798 82294 365854 82350
rect 365922 82294 365978 82350
rect 365798 82170 365854 82226
rect 365922 82170 365978 82226
rect 365798 82046 365854 82102
rect 365922 82046 365978 82102
rect 365798 81922 365854 81978
rect 365922 81922 365978 81978
rect 396518 82294 396574 82350
rect 396642 82294 396698 82350
rect 396518 82170 396574 82226
rect 396642 82170 396698 82226
rect 396518 82046 396574 82102
rect 396642 82046 396698 82102
rect 396518 81922 396574 81978
rect 396642 81922 396698 81978
rect 427238 82294 427294 82350
rect 427362 82294 427418 82350
rect 427238 82170 427294 82226
rect 427362 82170 427418 82226
rect 427238 82046 427294 82102
rect 427362 82046 427418 82102
rect 427238 81922 427294 81978
rect 427362 81922 427418 81978
rect 457958 82294 458014 82350
rect 458082 82294 458138 82350
rect 457958 82170 458014 82226
rect 458082 82170 458138 82226
rect 457958 82046 458014 82102
rect 458082 82046 458138 82102
rect 457958 81922 458014 81978
rect 458082 81922 458138 81978
rect 488678 82294 488734 82350
rect 488802 82294 488858 82350
rect 488678 82170 488734 82226
rect 488802 82170 488858 82226
rect 488678 82046 488734 82102
rect 488802 82046 488858 82102
rect 488678 81922 488734 81978
rect 488802 81922 488858 81978
rect 519398 82294 519454 82350
rect 519522 82294 519578 82350
rect 519398 82170 519454 82226
rect 519522 82170 519578 82226
rect 519398 82046 519454 82102
rect 519522 82046 519578 82102
rect 519398 81922 519454 81978
rect 519522 81922 519578 81978
rect 550118 82294 550174 82350
rect 550242 82294 550298 82350
rect 550118 82170 550174 82226
rect 550242 82170 550298 82226
rect 550118 82046 550174 82102
rect 550242 82046 550298 82102
rect 550118 81922 550174 81978
rect 550242 81922 550298 81978
rect 5514 76294 5570 76350
rect 5638 76294 5694 76350
rect 5762 76294 5818 76350
rect 5886 76294 5942 76350
rect 5514 76170 5570 76226
rect 5638 76170 5694 76226
rect 5762 76170 5818 76226
rect 5886 76170 5942 76226
rect 5514 76046 5570 76102
rect 5638 76046 5694 76102
rect 5762 76046 5818 76102
rect 5886 76046 5942 76102
rect 5514 75922 5570 75978
rect 5638 75922 5694 75978
rect 5762 75922 5818 75978
rect 5886 75922 5942 75978
rect -860 58294 -804 58350
rect -736 58294 -680 58350
rect -612 58294 -556 58350
rect -488 58294 -432 58350
rect -860 58170 -804 58226
rect -736 58170 -680 58226
rect -612 58170 -556 58226
rect -488 58170 -432 58226
rect -860 58046 -804 58102
rect -736 58046 -680 58102
rect -612 58046 -556 58102
rect -488 58046 -432 58102
rect -860 57922 -804 57978
rect -736 57922 -680 57978
rect -612 57922 -556 57978
rect -488 57922 -432 57978
rect 12518 76294 12574 76350
rect 12642 76294 12698 76350
rect 12518 76170 12574 76226
rect 12642 76170 12698 76226
rect 12518 76046 12574 76102
rect 12642 76046 12698 76102
rect 12518 75922 12574 75978
rect 12642 75922 12698 75978
rect 43238 76294 43294 76350
rect 43362 76294 43418 76350
rect 43238 76170 43294 76226
rect 43362 76170 43418 76226
rect 43238 76046 43294 76102
rect 43362 76046 43418 76102
rect 43238 75922 43294 75978
rect 43362 75922 43418 75978
rect 73958 76294 74014 76350
rect 74082 76294 74138 76350
rect 73958 76170 74014 76226
rect 74082 76170 74138 76226
rect 73958 76046 74014 76102
rect 74082 76046 74138 76102
rect 73958 75922 74014 75978
rect 74082 75922 74138 75978
rect 104678 76294 104734 76350
rect 104802 76294 104858 76350
rect 104678 76170 104734 76226
rect 104802 76170 104858 76226
rect 104678 76046 104734 76102
rect 104802 76046 104858 76102
rect 104678 75922 104734 75978
rect 104802 75922 104858 75978
rect 135398 76294 135454 76350
rect 135522 76294 135578 76350
rect 135398 76170 135454 76226
rect 135522 76170 135578 76226
rect 135398 76046 135454 76102
rect 135522 76046 135578 76102
rect 135398 75922 135454 75978
rect 135522 75922 135578 75978
rect 166118 76294 166174 76350
rect 166242 76294 166298 76350
rect 166118 76170 166174 76226
rect 166242 76170 166298 76226
rect 166118 76046 166174 76102
rect 166242 76046 166298 76102
rect 166118 75922 166174 75978
rect 166242 75922 166298 75978
rect 196838 76294 196894 76350
rect 196962 76294 197018 76350
rect 196838 76170 196894 76226
rect 196962 76170 197018 76226
rect 196838 76046 196894 76102
rect 196962 76046 197018 76102
rect 196838 75922 196894 75978
rect 196962 75922 197018 75978
rect 227558 76294 227614 76350
rect 227682 76294 227738 76350
rect 227558 76170 227614 76226
rect 227682 76170 227738 76226
rect 227558 76046 227614 76102
rect 227682 76046 227738 76102
rect 227558 75922 227614 75978
rect 227682 75922 227738 75978
rect 258278 76294 258334 76350
rect 258402 76294 258458 76350
rect 258278 76170 258334 76226
rect 258402 76170 258458 76226
rect 258278 76046 258334 76102
rect 258402 76046 258458 76102
rect 258278 75922 258334 75978
rect 258402 75922 258458 75978
rect 288998 76294 289054 76350
rect 289122 76294 289178 76350
rect 288998 76170 289054 76226
rect 289122 76170 289178 76226
rect 288998 76046 289054 76102
rect 289122 76046 289178 76102
rect 288998 75922 289054 75978
rect 289122 75922 289178 75978
rect 319718 76294 319774 76350
rect 319842 76294 319898 76350
rect 319718 76170 319774 76226
rect 319842 76170 319898 76226
rect 319718 76046 319774 76102
rect 319842 76046 319898 76102
rect 319718 75922 319774 75978
rect 319842 75922 319898 75978
rect 350438 76294 350494 76350
rect 350562 76294 350618 76350
rect 350438 76170 350494 76226
rect 350562 76170 350618 76226
rect 350438 76046 350494 76102
rect 350562 76046 350618 76102
rect 350438 75922 350494 75978
rect 350562 75922 350618 75978
rect 381158 76294 381214 76350
rect 381282 76294 381338 76350
rect 381158 76170 381214 76226
rect 381282 76170 381338 76226
rect 381158 76046 381214 76102
rect 381282 76046 381338 76102
rect 381158 75922 381214 75978
rect 381282 75922 381338 75978
rect 411878 76294 411934 76350
rect 412002 76294 412058 76350
rect 411878 76170 411934 76226
rect 412002 76170 412058 76226
rect 411878 76046 411934 76102
rect 412002 76046 412058 76102
rect 411878 75922 411934 75978
rect 412002 75922 412058 75978
rect 442598 76294 442654 76350
rect 442722 76294 442778 76350
rect 442598 76170 442654 76226
rect 442722 76170 442778 76226
rect 442598 76046 442654 76102
rect 442722 76046 442778 76102
rect 442598 75922 442654 75978
rect 442722 75922 442778 75978
rect 473318 76294 473374 76350
rect 473442 76294 473498 76350
rect 473318 76170 473374 76226
rect 473442 76170 473498 76226
rect 473318 76046 473374 76102
rect 473442 76046 473498 76102
rect 473318 75922 473374 75978
rect 473442 75922 473498 75978
rect 504038 76294 504094 76350
rect 504162 76294 504218 76350
rect 504038 76170 504094 76226
rect 504162 76170 504218 76226
rect 504038 76046 504094 76102
rect 504162 76046 504218 76102
rect 504038 75922 504094 75978
rect 504162 75922 504218 75978
rect 534758 76294 534814 76350
rect 534882 76294 534938 76350
rect 534758 76170 534814 76226
rect 534882 76170 534938 76226
rect 534758 76046 534814 76102
rect 534882 76046 534938 76102
rect 534758 75922 534814 75978
rect 534882 75922 534938 75978
rect 565478 76294 565534 76350
rect 565602 76294 565658 76350
rect 565478 76170 565534 76226
rect 565602 76170 565658 76226
rect 565478 76046 565534 76102
rect 565602 76046 565658 76102
rect 565478 75922 565534 75978
rect 565602 75922 565658 75978
rect 592914 100294 592970 100350
rect 593038 100294 593094 100350
rect 593162 100294 593218 100350
rect 593286 100294 593342 100350
rect 592914 100170 592970 100226
rect 593038 100170 593094 100226
rect 593162 100170 593218 100226
rect 593286 100170 593342 100226
rect 592914 100046 592970 100102
rect 593038 100046 593094 100102
rect 593162 100046 593218 100102
rect 593286 100046 593342 100102
rect 592914 99922 592970 99978
rect 593038 99922 593094 99978
rect 593162 99922 593218 99978
rect 593286 99922 593342 99978
rect 592914 82294 592970 82350
rect 593038 82294 593094 82350
rect 593162 82294 593218 82350
rect 593286 82294 593342 82350
rect 592914 82170 592970 82226
rect 593038 82170 593094 82226
rect 593162 82170 593218 82226
rect 593286 82170 593342 82226
rect 592914 82046 592970 82102
rect 593038 82046 593094 82102
rect 593162 82046 593218 82102
rect 593286 82046 593342 82102
rect 592914 81922 592970 81978
rect 593038 81922 593094 81978
rect 593162 81922 593218 81978
rect 593286 81922 593342 81978
rect 589194 76294 589250 76350
rect 589318 76294 589374 76350
rect 589442 76294 589498 76350
rect 589566 76294 589622 76350
rect 589194 76170 589250 76226
rect 589318 76170 589374 76226
rect 589442 76170 589498 76226
rect 589566 76170 589622 76226
rect 589194 76046 589250 76102
rect 589318 76046 589374 76102
rect 589442 76046 589498 76102
rect 589566 76046 589622 76102
rect 589194 75922 589250 75978
rect 589318 75922 589374 75978
rect 589442 75922 589498 75978
rect 589566 75922 589622 75978
rect 27878 64294 27934 64350
rect 28002 64294 28058 64350
rect 27878 64170 27934 64226
rect 28002 64170 28058 64226
rect 27878 64046 27934 64102
rect 28002 64046 28058 64102
rect 27878 63922 27934 63978
rect 28002 63922 28058 63978
rect 58598 64294 58654 64350
rect 58722 64294 58778 64350
rect 58598 64170 58654 64226
rect 58722 64170 58778 64226
rect 58598 64046 58654 64102
rect 58722 64046 58778 64102
rect 58598 63922 58654 63978
rect 58722 63922 58778 63978
rect 89318 64294 89374 64350
rect 89442 64294 89498 64350
rect 89318 64170 89374 64226
rect 89442 64170 89498 64226
rect 89318 64046 89374 64102
rect 89442 64046 89498 64102
rect 89318 63922 89374 63978
rect 89442 63922 89498 63978
rect 120038 64294 120094 64350
rect 120162 64294 120218 64350
rect 120038 64170 120094 64226
rect 120162 64170 120218 64226
rect 120038 64046 120094 64102
rect 120162 64046 120218 64102
rect 120038 63922 120094 63978
rect 120162 63922 120218 63978
rect 150758 64294 150814 64350
rect 150882 64294 150938 64350
rect 150758 64170 150814 64226
rect 150882 64170 150938 64226
rect 150758 64046 150814 64102
rect 150882 64046 150938 64102
rect 150758 63922 150814 63978
rect 150882 63922 150938 63978
rect 181478 64294 181534 64350
rect 181602 64294 181658 64350
rect 181478 64170 181534 64226
rect 181602 64170 181658 64226
rect 181478 64046 181534 64102
rect 181602 64046 181658 64102
rect 181478 63922 181534 63978
rect 181602 63922 181658 63978
rect 212198 64294 212254 64350
rect 212322 64294 212378 64350
rect 212198 64170 212254 64226
rect 212322 64170 212378 64226
rect 212198 64046 212254 64102
rect 212322 64046 212378 64102
rect 212198 63922 212254 63978
rect 212322 63922 212378 63978
rect 242918 64294 242974 64350
rect 243042 64294 243098 64350
rect 242918 64170 242974 64226
rect 243042 64170 243098 64226
rect 242918 64046 242974 64102
rect 243042 64046 243098 64102
rect 242918 63922 242974 63978
rect 243042 63922 243098 63978
rect 273638 64294 273694 64350
rect 273762 64294 273818 64350
rect 273638 64170 273694 64226
rect 273762 64170 273818 64226
rect 273638 64046 273694 64102
rect 273762 64046 273818 64102
rect 273638 63922 273694 63978
rect 273762 63922 273818 63978
rect 304358 64294 304414 64350
rect 304482 64294 304538 64350
rect 304358 64170 304414 64226
rect 304482 64170 304538 64226
rect 304358 64046 304414 64102
rect 304482 64046 304538 64102
rect 304358 63922 304414 63978
rect 304482 63922 304538 63978
rect 335078 64294 335134 64350
rect 335202 64294 335258 64350
rect 335078 64170 335134 64226
rect 335202 64170 335258 64226
rect 335078 64046 335134 64102
rect 335202 64046 335258 64102
rect 335078 63922 335134 63978
rect 335202 63922 335258 63978
rect 365798 64294 365854 64350
rect 365922 64294 365978 64350
rect 365798 64170 365854 64226
rect 365922 64170 365978 64226
rect 365798 64046 365854 64102
rect 365922 64046 365978 64102
rect 365798 63922 365854 63978
rect 365922 63922 365978 63978
rect 396518 64294 396574 64350
rect 396642 64294 396698 64350
rect 396518 64170 396574 64226
rect 396642 64170 396698 64226
rect 396518 64046 396574 64102
rect 396642 64046 396698 64102
rect 396518 63922 396574 63978
rect 396642 63922 396698 63978
rect 427238 64294 427294 64350
rect 427362 64294 427418 64350
rect 427238 64170 427294 64226
rect 427362 64170 427418 64226
rect 427238 64046 427294 64102
rect 427362 64046 427418 64102
rect 427238 63922 427294 63978
rect 427362 63922 427418 63978
rect 457958 64294 458014 64350
rect 458082 64294 458138 64350
rect 457958 64170 458014 64226
rect 458082 64170 458138 64226
rect 457958 64046 458014 64102
rect 458082 64046 458138 64102
rect 457958 63922 458014 63978
rect 458082 63922 458138 63978
rect 488678 64294 488734 64350
rect 488802 64294 488858 64350
rect 488678 64170 488734 64226
rect 488802 64170 488858 64226
rect 488678 64046 488734 64102
rect 488802 64046 488858 64102
rect 488678 63922 488734 63978
rect 488802 63922 488858 63978
rect 519398 64294 519454 64350
rect 519522 64294 519578 64350
rect 519398 64170 519454 64226
rect 519522 64170 519578 64226
rect 519398 64046 519454 64102
rect 519522 64046 519578 64102
rect 519398 63922 519454 63978
rect 519522 63922 519578 63978
rect 550118 64294 550174 64350
rect 550242 64294 550298 64350
rect 550118 64170 550174 64226
rect 550242 64170 550298 64226
rect 550118 64046 550174 64102
rect 550242 64046 550298 64102
rect 550118 63922 550174 63978
rect 550242 63922 550298 63978
rect 5514 58294 5570 58350
rect 5638 58294 5694 58350
rect 5762 58294 5818 58350
rect 5886 58294 5942 58350
rect 5514 58170 5570 58226
rect 5638 58170 5694 58226
rect 5762 58170 5818 58226
rect 5886 58170 5942 58226
rect 5514 58046 5570 58102
rect 5638 58046 5694 58102
rect 5762 58046 5818 58102
rect 5886 58046 5942 58102
rect 5514 57922 5570 57978
rect 5638 57922 5694 57978
rect 5762 57922 5818 57978
rect 5886 57922 5942 57978
rect -860 40294 -804 40350
rect -736 40294 -680 40350
rect -612 40294 -556 40350
rect -488 40294 -432 40350
rect -860 40170 -804 40226
rect -736 40170 -680 40226
rect -612 40170 -556 40226
rect -488 40170 -432 40226
rect -860 40046 -804 40102
rect -736 40046 -680 40102
rect -612 40046 -556 40102
rect -488 40046 -432 40102
rect -860 39922 -804 39978
rect -736 39922 -680 39978
rect -612 39922 -556 39978
rect -488 39922 -432 39978
rect 12518 58294 12574 58350
rect 12642 58294 12698 58350
rect 12518 58170 12574 58226
rect 12642 58170 12698 58226
rect 12518 58046 12574 58102
rect 12642 58046 12698 58102
rect 12518 57922 12574 57978
rect 12642 57922 12698 57978
rect 43238 58294 43294 58350
rect 43362 58294 43418 58350
rect 43238 58170 43294 58226
rect 43362 58170 43418 58226
rect 43238 58046 43294 58102
rect 43362 58046 43418 58102
rect 43238 57922 43294 57978
rect 43362 57922 43418 57978
rect 73958 58294 74014 58350
rect 74082 58294 74138 58350
rect 73958 58170 74014 58226
rect 74082 58170 74138 58226
rect 73958 58046 74014 58102
rect 74082 58046 74138 58102
rect 73958 57922 74014 57978
rect 74082 57922 74138 57978
rect 104678 58294 104734 58350
rect 104802 58294 104858 58350
rect 104678 58170 104734 58226
rect 104802 58170 104858 58226
rect 104678 58046 104734 58102
rect 104802 58046 104858 58102
rect 104678 57922 104734 57978
rect 104802 57922 104858 57978
rect 135398 58294 135454 58350
rect 135522 58294 135578 58350
rect 135398 58170 135454 58226
rect 135522 58170 135578 58226
rect 135398 58046 135454 58102
rect 135522 58046 135578 58102
rect 135398 57922 135454 57978
rect 135522 57922 135578 57978
rect 166118 58294 166174 58350
rect 166242 58294 166298 58350
rect 166118 58170 166174 58226
rect 166242 58170 166298 58226
rect 166118 58046 166174 58102
rect 166242 58046 166298 58102
rect 166118 57922 166174 57978
rect 166242 57922 166298 57978
rect 196838 58294 196894 58350
rect 196962 58294 197018 58350
rect 196838 58170 196894 58226
rect 196962 58170 197018 58226
rect 196838 58046 196894 58102
rect 196962 58046 197018 58102
rect 196838 57922 196894 57978
rect 196962 57922 197018 57978
rect 227558 58294 227614 58350
rect 227682 58294 227738 58350
rect 227558 58170 227614 58226
rect 227682 58170 227738 58226
rect 227558 58046 227614 58102
rect 227682 58046 227738 58102
rect 227558 57922 227614 57978
rect 227682 57922 227738 57978
rect 258278 58294 258334 58350
rect 258402 58294 258458 58350
rect 258278 58170 258334 58226
rect 258402 58170 258458 58226
rect 258278 58046 258334 58102
rect 258402 58046 258458 58102
rect 258278 57922 258334 57978
rect 258402 57922 258458 57978
rect 288998 58294 289054 58350
rect 289122 58294 289178 58350
rect 288998 58170 289054 58226
rect 289122 58170 289178 58226
rect 288998 58046 289054 58102
rect 289122 58046 289178 58102
rect 288998 57922 289054 57978
rect 289122 57922 289178 57978
rect 319718 58294 319774 58350
rect 319842 58294 319898 58350
rect 319718 58170 319774 58226
rect 319842 58170 319898 58226
rect 319718 58046 319774 58102
rect 319842 58046 319898 58102
rect 319718 57922 319774 57978
rect 319842 57922 319898 57978
rect 350438 58294 350494 58350
rect 350562 58294 350618 58350
rect 350438 58170 350494 58226
rect 350562 58170 350618 58226
rect 350438 58046 350494 58102
rect 350562 58046 350618 58102
rect 350438 57922 350494 57978
rect 350562 57922 350618 57978
rect 381158 58294 381214 58350
rect 381282 58294 381338 58350
rect 381158 58170 381214 58226
rect 381282 58170 381338 58226
rect 381158 58046 381214 58102
rect 381282 58046 381338 58102
rect 381158 57922 381214 57978
rect 381282 57922 381338 57978
rect 411878 58294 411934 58350
rect 412002 58294 412058 58350
rect 411878 58170 411934 58226
rect 412002 58170 412058 58226
rect 411878 58046 411934 58102
rect 412002 58046 412058 58102
rect 411878 57922 411934 57978
rect 412002 57922 412058 57978
rect 442598 58294 442654 58350
rect 442722 58294 442778 58350
rect 442598 58170 442654 58226
rect 442722 58170 442778 58226
rect 442598 58046 442654 58102
rect 442722 58046 442778 58102
rect 442598 57922 442654 57978
rect 442722 57922 442778 57978
rect 473318 58294 473374 58350
rect 473442 58294 473498 58350
rect 473318 58170 473374 58226
rect 473442 58170 473498 58226
rect 473318 58046 473374 58102
rect 473442 58046 473498 58102
rect 473318 57922 473374 57978
rect 473442 57922 473498 57978
rect 504038 58294 504094 58350
rect 504162 58294 504218 58350
rect 504038 58170 504094 58226
rect 504162 58170 504218 58226
rect 504038 58046 504094 58102
rect 504162 58046 504218 58102
rect 504038 57922 504094 57978
rect 504162 57922 504218 57978
rect 534758 58294 534814 58350
rect 534882 58294 534938 58350
rect 534758 58170 534814 58226
rect 534882 58170 534938 58226
rect 534758 58046 534814 58102
rect 534882 58046 534938 58102
rect 534758 57922 534814 57978
rect 534882 57922 534938 57978
rect 565478 58294 565534 58350
rect 565602 58294 565658 58350
rect 565478 58170 565534 58226
rect 565602 58170 565658 58226
rect 565478 58046 565534 58102
rect 565602 58046 565658 58102
rect 565478 57922 565534 57978
rect 565602 57922 565658 57978
rect 589194 58294 589250 58350
rect 589318 58294 589374 58350
rect 589442 58294 589498 58350
rect 589566 58294 589622 58350
rect 589194 58170 589250 58226
rect 589318 58170 589374 58226
rect 589442 58170 589498 58226
rect 589566 58170 589622 58226
rect 589194 58046 589250 58102
rect 589318 58046 589374 58102
rect 589442 58046 589498 58102
rect 589566 58046 589622 58102
rect 589194 57922 589250 57978
rect 589318 57922 589374 57978
rect 589442 57922 589498 57978
rect 589566 57922 589622 57978
rect 27878 46294 27934 46350
rect 28002 46294 28058 46350
rect 27878 46170 27934 46226
rect 28002 46170 28058 46226
rect 27878 46046 27934 46102
rect 28002 46046 28058 46102
rect 27878 45922 27934 45978
rect 28002 45922 28058 45978
rect 58598 46294 58654 46350
rect 58722 46294 58778 46350
rect 58598 46170 58654 46226
rect 58722 46170 58778 46226
rect 58598 46046 58654 46102
rect 58722 46046 58778 46102
rect 58598 45922 58654 45978
rect 58722 45922 58778 45978
rect 89318 46294 89374 46350
rect 89442 46294 89498 46350
rect 89318 46170 89374 46226
rect 89442 46170 89498 46226
rect 89318 46046 89374 46102
rect 89442 46046 89498 46102
rect 89318 45922 89374 45978
rect 89442 45922 89498 45978
rect 120038 46294 120094 46350
rect 120162 46294 120218 46350
rect 120038 46170 120094 46226
rect 120162 46170 120218 46226
rect 120038 46046 120094 46102
rect 120162 46046 120218 46102
rect 120038 45922 120094 45978
rect 120162 45922 120218 45978
rect 150758 46294 150814 46350
rect 150882 46294 150938 46350
rect 150758 46170 150814 46226
rect 150882 46170 150938 46226
rect 150758 46046 150814 46102
rect 150882 46046 150938 46102
rect 150758 45922 150814 45978
rect 150882 45922 150938 45978
rect 181478 46294 181534 46350
rect 181602 46294 181658 46350
rect 181478 46170 181534 46226
rect 181602 46170 181658 46226
rect 181478 46046 181534 46102
rect 181602 46046 181658 46102
rect 181478 45922 181534 45978
rect 181602 45922 181658 45978
rect 212198 46294 212254 46350
rect 212322 46294 212378 46350
rect 212198 46170 212254 46226
rect 212322 46170 212378 46226
rect 212198 46046 212254 46102
rect 212322 46046 212378 46102
rect 212198 45922 212254 45978
rect 212322 45922 212378 45978
rect 242918 46294 242974 46350
rect 243042 46294 243098 46350
rect 242918 46170 242974 46226
rect 243042 46170 243098 46226
rect 242918 46046 242974 46102
rect 243042 46046 243098 46102
rect 242918 45922 242974 45978
rect 243042 45922 243098 45978
rect 273638 46294 273694 46350
rect 273762 46294 273818 46350
rect 273638 46170 273694 46226
rect 273762 46170 273818 46226
rect 273638 46046 273694 46102
rect 273762 46046 273818 46102
rect 273638 45922 273694 45978
rect 273762 45922 273818 45978
rect 304358 46294 304414 46350
rect 304482 46294 304538 46350
rect 304358 46170 304414 46226
rect 304482 46170 304538 46226
rect 304358 46046 304414 46102
rect 304482 46046 304538 46102
rect 304358 45922 304414 45978
rect 304482 45922 304538 45978
rect 335078 46294 335134 46350
rect 335202 46294 335258 46350
rect 335078 46170 335134 46226
rect 335202 46170 335258 46226
rect 335078 46046 335134 46102
rect 335202 46046 335258 46102
rect 335078 45922 335134 45978
rect 335202 45922 335258 45978
rect 365798 46294 365854 46350
rect 365922 46294 365978 46350
rect 365798 46170 365854 46226
rect 365922 46170 365978 46226
rect 365798 46046 365854 46102
rect 365922 46046 365978 46102
rect 365798 45922 365854 45978
rect 365922 45922 365978 45978
rect 396518 46294 396574 46350
rect 396642 46294 396698 46350
rect 396518 46170 396574 46226
rect 396642 46170 396698 46226
rect 396518 46046 396574 46102
rect 396642 46046 396698 46102
rect 396518 45922 396574 45978
rect 396642 45922 396698 45978
rect 427238 46294 427294 46350
rect 427362 46294 427418 46350
rect 427238 46170 427294 46226
rect 427362 46170 427418 46226
rect 427238 46046 427294 46102
rect 427362 46046 427418 46102
rect 427238 45922 427294 45978
rect 427362 45922 427418 45978
rect 457958 46294 458014 46350
rect 458082 46294 458138 46350
rect 457958 46170 458014 46226
rect 458082 46170 458138 46226
rect 457958 46046 458014 46102
rect 458082 46046 458138 46102
rect 457958 45922 458014 45978
rect 458082 45922 458138 45978
rect 488678 46294 488734 46350
rect 488802 46294 488858 46350
rect 488678 46170 488734 46226
rect 488802 46170 488858 46226
rect 488678 46046 488734 46102
rect 488802 46046 488858 46102
rect 488678 45922 488734 45978
rect 488802 45922 488858 45978
rect 519398 46294 519454 46350
rect 519522 46294 519578 46350
rect 519398 46170 519454 46226
rect 519522 46170 519578 46226
rect 519398 46046 519454 46102
rect 519522 46046 519578 46102
rect 519398 45922 519454 45978
rect 519522 45922 519578 45978
rect 550118 46294 550174 46350
rect 550242 46294 550298 46350
rect 550118 46170 550174 46226
rect 550242 46170 550298 46226
rect 550118 46046 550174 46102
rect 550242 46046 550298 46102
rect 550118 45922 550174 45978
rect 550242 45922 550298 45978
rect 5514 40294 5570 40350
rect 5638 40294 5694 40350
rect 5762 40294 5818 40350
rect 5886 40294 5942 40350
rect 5514 40170 5570 40226
rect 5638 40170 5694 40226
rect 5762 40170 5818 40226
rect 5886 40170 5942 40226
rect 5514 40046 5570 40102
rect 5638 40046 5694 40102
rect 5762 40046 5818 40102
rect 5886 40046 5942 40102
rect 5514 39922 5570 39978
rect 5638 39922 5694 39978
rect 5762 39922 5818 39978
rect 5886 39922 5942 39978
rect -860 22294 -804 22350
rect -736 22294 -680 22350
rect -612 22294 -556 22350
rect -488 22294 -432 22350
rect -860 22170 -804 22226
rect -736 22170 -680 22226
rect -612 22170 -556 22226
rect -488 22170 -432 22226
rect -860 22046 -804 22102
rect -736 22046 -680 22102
rect -612 22046 -556 22102
rect -488 22046 -432 22102
rect -860 21922 -804 21978
rect -736 21922 -680 21978
rect -612 21922 -556 21978
rect -488 21922 -432 21978
rect -860 4294 -804 4350
rect -736 4294 -680 4350
rect -612 4294 -556 4350
rect -488 4294 -432 4350
rect -860 4170 -804 4226
rect -736 4170 -680 4226
rect -612 4170 -556 4226
rect -488 4170 -432 4226
rect -860 4046 -804 4102
rect -736 4046 -680 4102
rect -612 4046 -556 4102
rect -488 4046 -432 4102
rect -860 3922 -804 3978
rect -736 3922 -680 3978
rect -612 3922 -556 3978
rect -488 3922 -432 3978
rect -860 -216 -804 -160
rect -736 -216 -680 -160
rect -612 -216 -556 -160
rect -488 -216 -432 -160
rect -860 -340 -804 -284
rect -736 -340 -680 -284
rect -612 -340 -556 -284
rect -488 -340 -432 -284
rect -860 -464 -804 -408
rect -736 -464 -680 -408
rect -612 -464 -556 -408
rect -488 -464 -432 -408
rect -860 -588 -804 -532
rect -736 -588 -680 -532
rect -612 -588 -556 -532
rect -488 -588 -432 -532
rect 12518 40294 12574 40350
rect 12642 40294 12698 40350
rect 12518 40170 12574 40226
rect 12642 40170 12698 40226
rect 12518 40046 12574 40102
rect 12642 40046 12698 40102
rect 12518 39922 12574 39978
rect 12642 39922 12698 39978
rect 43238 40294 43294 40350
rect 43362 40294 43418 40350
rect 43238 40170 43294 40226
rect 43362 40170 43418 40226
rect 43238 40046 43294 40102
rect 43362 40046 43418 40102
rect 43238 39922 43294 39978
rect 43362 39922 43418 39978
rect 73958 40294 74014 40350
rect 74082 40294 74138 40350
rect 73958 40170 74014 40226
rect 74082 40170 74138 40226
rect 73958 40046 74014 40102
rect 74082 40046 74138 40102
rect 73958 39922 74014 39978
rect 74082 39922 74138 39978
rect 104678 40294 104734 40350
rect 104802 40294 104858 40350
rect 104678 40170 104734 40226
rect 104802 40170 104858 40226
rect 104678 40046 104734 40102
rect 104802 40046 104858 40102
rect 104678 39922 104734 39978
rect 104802 39922 104858 39978
rect 135398 40294 135454 40350
rect 135522 40294 135578 40350
rect 135398 40170 135454 40226
rect 135522 40170 135578 40226
rect 135398 40046 135454 40102
rect 135522 40046 135578 40102
rect 135398 39922 135454 39978
rect 135522 39922 135578 39978
rect 166118 40294 166174 40350
rect 166242 40294 166298 40350
rect 166118 40170 166174 40226
rect 166242 40170 166298 40226
rect 166118 40046 166174 40102
rect 166242 40046 166298 40102
rect 166118 39922 166174 39978
rect 166242 39922 166298 39978
rect 196838 40294 196894 40350
rect 196962 40294 197018 40350
rect 196838 40170 196894 40226
rect 196962 40170 197018 40226
rect 196838 40046 196894 40102
rect 196962 40046 197018 40102
rect 196838 39922 196894 39978
rect 196962 39922 197018 39978
rect 227558 40294 227614 40350
rect 227682 40294 227738 40350
rect 227558 40170 227614 40226
rect 227682 40170 227738 40226
rect 227558 40046 227614 40102
rect 227682 40046 227738 40102
rect 227558 39922 227614 39978
rect 227682 39922 227738 39978
rect 258278 40294 258334 40350
rect 258402 40294 258458 40350
rect 258278 40170 258334 40226
rect 258402 40170 258458 40226
rect 258278 40046 258334 40102
rect 258402 40046 258458 40102
rect 258278 39922 258334 39978
rect 258402 39922 258458 39978
rect 288998 40294 289054 40350
rect 289122 40294 289178 40350
rect 288998 40170 289054 40226
rect 289122 40170 289178 40226
rect 288998 40046 289054 40102
rect 289122 40046 289178 40102
rect 288998 39922 289054 39978
rect 289122 39922 289178 39978
rect 319718 40294 319774 40350
rect 319842 40294 319898 40350
rect 319718 40170 319774 40226
rect 319842 40170 319898 40226
rect 319718 40046 319774 40102
rect 319842 40046 319898 40102
rect 319718 39922 319774 39978
rect 319842 39922 319898 39978
rect 350438 40294 350494 40350
rect 350562 40294 350618 40350
rect 350438 40170 350494 40226
rect 350562 40170 350618 40226
rect 350438 40046 350494 40102
rect 350562 40046 350618 40102
rect 350438 39922 350494 39978
rect 350562 39922 350618 39978
rect 381158 40294 381214 40350
rect 381282 40294 381338 40350
rect 381158 40170 381214 40226
rect 381282 40170 381338 40226
rect 381158 40046 381214 40102
rect 381282 40046 381338 40102
rect 381158 39922 381214 39978
rect 381282 39922 381338 39978
rect 411878 40294 411934 40350
rect 412002 40294 412058 40350
rect 411878 40170 411934 40226
rect 412002 40170 412058 40226
rect 411878 40046 411934 40102
rect 412002 40046 412058 40102
rect 411878 39922 411934 39978
rect 412002 39922 412058 39978
rect 442598 40294 442654 40350
rect 442722 40294 442778 40350
rect 442598 40170 442654 40226
rect 442722 40170 442778 40226
rect 442598 40046 442654 40102
rect 442722 40046 442778 40102
rect 442598 39922 442654 39978
rect 442722 39922 442778 39978
rect 473318 40294 473374 40350
rect 473442 40294 473498 40350
rect 473318 40170 473374 40226
rect 473442 40170 473498 40226
rect 473318 40046 473374 40102
rect 473442 40046 473498 40102
rect 473318 39922 473374 39978
rect 473442 39922 473498 39978
rect 504038 40294 504094 40350
rect 504162 40294 504218 40350
rect 504038 40170 504094 40226
rect 504162 40170 504218 40226
rect 504038 40046 504094 40102
rect 504162 40046 504218 40102
rect 504038 39922 504094 39978
rect 504162 39922 504218 39978
rect 534758 40294 534814 40350
rect 534882 40294 534938 40350
rect 534758 40170 534814 40226
rect 534882 40170 534938 40226
rect 534758 40046 534814 40102
rect 534882 40046 534938 40102
rect 534758 39922 534814 39978
rect 534882 39922 534938 39978
rect 565478 40294 565534 40350
rect 565602 40294 565658 40350
rect 565478 40170 565534 40226
rect 565602 40170 565658 40226
rect 565478 40046 565534 40102
rect 565602 40046 565658 40102
rect 565478 39922 565534 39978
rect 565602 39922 565658 39978
rect 592914 64294 592970 64350
rect 593038 64294 593094 64350
rect 593162 64294 593218 64350
rect 593286 64294 593342 64350
rect 592914 64170 592970 64226
rect 593038 64170 593094 64226
rect 593162 64170 593218 64226
rect 593286 64170 593342 64226
rect 592914 64046 592970 64102
rect 593038 64046 593094 64102
rect 593162 64046 593218 64102
rect 593286 64046 593342 64102
rect 592914 63922 592970 63978
rect 593038 63922 593094 63978
rect 593162 63922 593218 63978
rect 593286 63922 593342 63978
rect 589194 40294 589250 40350
rect 589318 40294 589374 40350
rect 589442 40294 589498 40350
rect 589566 40294 589622 40350
rect 589194 40170 589250 40226
rect 589318 40170 589374 40226
rect 589442 40170 589498 40226
rect 589566 40170 589622 40226
rect 589194 40046 589250 40102
rect 589318 40046 589374 40102
rect 589442 40046 589498 40102
rect 589566 40046 589622 40102
rect 589194 39922 589250 39978
rect 589318 39922 589374 39978
rect 589442 39922 589498 39978
rect 589566 39922 589622 39978
rect 27878 28294 27934 28350
rect 28002 28294 28058 28350
rect 27878 28170 27934 28226
rect 28002 28170 28058 28226
rect 27878 28046 27934 28102
rect 28002 28046 28058 28102
rect 27878 27922 27934 27978
rect 28002 27922 28058 27978
rect 58598 28294 58654 28350
rect 58722 28294 58778 28350
rect 58598 28170 58654 28226
rect 58722 28170 58778 28226
rect 58598 28046 58654 28102
rect 58722 28046 58778 28102
rect 58598 27922 58654 27978
rect 58722 27922 58778 27978
rect 89318 28294 89374 28350
rect 89442 28294 89498 28350
rect 89318 28170 89374 28226
rect 89442 28170 89498 28226
rect 89318 28046 89374 28102
rect 89442 28046 89498 28102
rect 89318 27922 89374 27978
rect 89442 27922 89498 27978
rect 120038 28294 120094 28350
rect 120162 28294 120218 28350
rect 120038 28170 120094 28226
rect 120162 28170 120218 28226
rect 120038 28046 120094 28102
rect 120162 28046 120218 28102
rect 120038 27922 120094 27978
rect 120162 27922 120218 27978
rect 150758 28294 150814 28350
rect 150882 28294 150938 28350
rect 150758 28170 150814 28226
rect 150882 28170 150938 28226
rect 150758 28046 150814 28102
rect 150882 28046 150938 28102
rect 150758 27922 150814 27978
rect 150882 27922 150938 27978
rect 181478 28294 181534 28350
rect 181602 28294 181658 28350
rect 181478 28170 181534 28226
rect 181602 28170 181658 28226
rect 181478 28046 181534 28102
rect 181602 28046 181658 28102
rect 181478 27922 181534 27978
rect 181602 27922 181658 27978
rect 212198 28294 212254 28350
rect 212322 28294 212378 28350
rect 212198 28170 212254 28226
rect 212322 28170 212378 28226
rect 212198 28046 212254 28102
rect 212322 28046 212378 28102
rect 212198 27922 212254 27978
rect 212322 27922 212378 27978
rect 242918 28294 242974 28350
rect 243042 28294 243098 28350
rect 242918 28170 242974 28226
rect 243042 28170 243098 28226
rect 242918 28046 242974 28102
rect 243042 28046 243098 28102
rect 242918 27922 242974 27978
rect 243042 27922 243098 27978
rect 273638 28294 273694 28350
rect 273762 28294 273818 28350
rect 273638 28170 273694 28226
rect 273762 28170 273818 28226
rect 273638 28046 273694 28102
rect 273762 28046 273818 28102
rect 273638 27922 273694 27978
rect 273762 27922 273818 27978
rect 304358 28294 304414 28350
rect 304482 28294 304538 28350
rect 304358 28170 304414 28226
rect 304482 28170 304538 28226
rect 304358 28046 304414 28102
rect 304482 28046 304538 28102
rect 304358 27922 304414 27978
rect 304482 27922 304538 27978
rect 335078 28294 335134 28350
rect 335202 28294 335258 28350
rect 335078 28170 335134 28226
rect 335202 28170 335258 28226
rect 335078 28046 335134 28102
rect 335202 28046 335258 28102
rect 335078 27922 335134 27978
rect 335202 27922 335258 27978
rect 365798 28294 365854 28350
rect 365922 28294 365978 28350
rect 365798 28170 365854 28226
rect 365922 28170 365978 28226
rect 365798 28046 365854 28102
rect 365922 28046 365978 28102
rect 365798 27922 365854 27978
rect 365922 27922 365978 27978
rect 396518 28294 396574 28350
rect 396642 28294 396698 28350
rect 396518 28170 396574 28226
rect 396642 28170 396698 28226
rect 396518 28046 396574 28102
rect 396642 28046 396698 28102
rect 396518 27922 396574 27978
rect 396642 27922 396698 27978
rect 427238 28294 427294 28350
rect 427362 28294 427418 28350
rect 427238 28170 427294 28226
rect 427362 28170 427418 28226
rect 427238 28046 427294 28102
rect 427362 28046 427418 28102
rect 427238 27922 427294 27978
rect 427362 27922 427418 27978
rect 457958 28294 458014 28350
rect 458082 28294 458138 28350
rect 457958 28170 458014 28226
rect 458082 28170 458138 28226
rect 457958 28046 458014 28102
rect 458082 28046 458138 28102
rect 457958 27922 458014 27978
rect 458082 27922 458138 27978
rect 488678 28294 488734 28350
rect 488802 28294 488858 28350
rect 488678 28170 488734 28226
rect 488802 28170 488858 28226
rect 488678 28046 488734 28102
rect 488802 28046 488858 28102
rect 488678 27922 488734 27978
rect 488802 27922 488858 27978
rect 519398 28294 519454 28350
rect 519522 28294 519578 28350
rect 519398 28170 519454 28226
rect 519522 28170 519578 28226
rect 519398 28046 519454 28102
rect 519522 28046 519578 28102
rect 519398 27922 519454 27978
rect 519522 27922 519578 27978
rect 550118 28294 550174 28350
rect 550242 28294 550298 28350
rect 550118 28170 550174 28226
rect 550242 28170 550298 28226
rect 550118 28046 550174 28102
rect 550242 28046 550298 28102
rect 550118 27922 550174 27978
rect 550242 27922 550298 27978
rect 5514 22294 5570 22350
rect 5638 22294 5694 22350
rect 5762 22294 5818 22350
rect 5886 22294 5942 22350
rect 5514 22170 5570 22226
rect 5638 22170 5694 22226
rect 5762 22170 5818 22226
rect 5886 22170 5942 22226
rect 5514 22046 5570 22102
rect 5638 22046 5694 22102
rect 5762 22046 5818 22102
rect 5886 22046 5942 22102
rect 5514 21922 5570 21978
rect 5638 21922 5694 21978
rect 5762 21922 5818 21978
rect 5886 21922 5942 21978
rect 12518 22294 12574 22350
rect 12642 22294 12698 22350
rect 12518 22170 12574 22226
rect 12642 22170 12698 22226
rect 12518 22046 12574 22102
rect 12642 22046 12698 22102
rect 12518 21922 12574 21978
rect 12642 21922 12698 21978
rect 43238 22294 43294 22350
rect 43362 22294 43418 22350
rect 43238 22170 43294 22226
rect 43362 22170 43418 22226
rect 43238 22046 43294 22102
rect 43362 22046 43418 22102
rect 43238 21922 43294 21978
rect 43362 21922 43418 21978
rect 73958 22294 74014 22350
rect 74082 22294 74138 22350
rect 73958 22170 74014 22226
rect 74082 22170 74138 22226
rect 73958 22046 74014 22102
rect 74082 22046 74138 22102
rect 73958 21922 74014 21978
rect 74082 21922 74138 21978
rect 104678 22294 104734 22350
rect 104802 22294 104858 22350
rect 104678 22170 104734 22226
rect 104802 22170 104858 22226
rect 104678 22046 104734 22102
rect 104802 22046 104858 22102
rect 104678 21922 104734 21978
rect 104802 21922 104858 21978
rect 135398 22294 135454 22350
rect 135522 22294 135578 22350
rect 135398 22170 135454 22226
rect 135522 22170 135578 22226
rect 135398 22046 135454 22102
rect 135522 22046 135578 22102
rect 135398 21922 135454 21978
rect 135522 21922 135578 21978
rect 166118 22294 166174 22350
rect 166242 22294 166298 22350
rect 166118 22170 166174 22226
rect 166242 22170 166298 22226
rect 166118 22046 166174 22102
rect 166242 22046 166298 22102
rect 166118 21922 166174 21978
rect 166242 21922 166298 21978
rect 196838 22294 196894 22350
rect 196962 22294 197018 22350
rect 196838 22170 196894 22226
rect 196962 22170 197018 22226
rect 196838 22046 196894 22102
rect 196962 22046 197018 22102
rect 196838 21922 196894 21978
rect 196962 21922 197018 21978
rect 227558 22294 227614 22350
rect 227682 22294 227738 22350
rect 227558 22170 227614 22226
rect 227682 22170 227738 22226
rect 227558 22046 227614 22102
rect 227682 22046 227738 22102
rect 227558 21922 227614 21978
rect 227682 21922 227738 21978
rect 258278 22294 258334 22350
rect 258402 22294 258458 22350
rect 258278 22170 258334 22226
rect 258402 22170 258458 22226
rect 258278 22046 258334 22102
rect 258402 22046 258458 22102
rect 258278 21922 258334 21978
rect 258402 21922 258458 21978
rect 288998 22294 289054 22350
rect 289122 22294 289178 22350
rect 288998 22170 289054 22226
rect 289122 22170 289178 22226
rect 288998 22046 289054 22102
rect 289122 22046 289178 22102
rect 288998 21922 289054 21978
rect 289122 21922 289178 21978
rect 319718 22294 319774 22350
rect 319842 22294 319898 22350
rect 319718 22170 319774 22226
rect 319842 22170 319898 22226
rect 319718 22046 319774 22102
rect 319842 22046 319898 22102
rect 319718 21922 319774 21978
rect 319842 21922 319898 21978
rect 350438 22294 350494 22350
rect 350562 22294 350618 22350
rect 350438 22170 350494 22226
rect 350562 22170 350618 22226
rect 350438 22046 350494 22102
rect 350562 22046 350618 22102
rect 350438 21922 350494 21978
rect 350562 21922 350618 21978
rect 381158 22294 381214 22350
rect 381282 22294 381338 22350
rect 381158 22170 381214 22226
rect 381282 22170 381338 22226
rect 381158 22046 381214 22102
rect 381282 22046 381338 22102
rect 381158 21922 381214 21978
rect 381282 21922 381338 21978
rect 411878 22294 411934 22350
rect 412002 22294 412058 22350
rect 411878 22170 411934 22226
rect 412002 22170 412058 22226
rect 411878 22046 411934 22102
rect 412002 22046 412058 22102
rect 411878 21922 411934 21978
rect 412002 21922 412058 21978
rect 442598 22294 442654 22350
rect 442722 22294 442778 22350
rect 442598 22170 442654 22226
rect 442722 22170 442778 22226
rect 442598 22046 442654 22102
rect 442722 22046 442778 22102
rect 442598 21922 442654 21978
rect 442722 21922 442778 21978
rect 473318 22294 473374 22350
rect 473442 22294 473498 22350
rect 473318 22170 473374 22226
rect 473442 22170 473498 22226
rect 473318 22046 473374 22102
rect 473442 22046 473498 22102
rect 473318 21922 473374 21978
rect 473442 21922 473498 21978
rect 504038 22294 504094 22350
rect 504162 22294 504218 22350
rect 504038 22170 504094 22226
rect 504162 22170 504218 22226
rect 504038 22046 504094 22102
rect 504162 22046 504218 22102
rect 504038 21922 504094 21978
rect 504162 21922 504218 21978
rect 534758 22294 534814 22350
rect 534882 22294 534938 22350
rect 534758 22170 534814 22226
rect 534882 22170 534938 22226
rect 534758 22046 534814 22102
rect 534882 22046 534938 22102
rect 534758 21922 534814 21978
rect 534882 21922 534938 21978
rect 565478 22294 565534 22350
rect 565602 22294 565658 22350
rect 565478 22170 565534 22226
rect 565602 22170 565658 22226
rect 565478 22046 565534 22102
rect 565602 22046 565658 22102
rect 565478 21922 565534 21978
rect 565602 21922 565658 21978
rect 589194 22294 589250 22350
rect 589318 22294 589374 22350
rect 589442 22294 589498 22350
rect 589566 22294 589622 22350
rect 589194 22170 589250 22226
rect 589318 22170 589374 22226
rect 589442 22170 589498 22226
rect 589566 22170 589622 22226
rect 589194 22046 589250 22102
rect 589318 22046 589374 22102
rect 589442 22046 589498 22102
rect 589566 22046 589622 22102
rect 589194 21922 589250 21978
rect 589318 21922 589374 21978
rect 589442 21922 589498 21978
rect 589566 21922 589622 21978
rect 5514 4294 5570 4350
rect 5638 4294 5694 4350
rect 5762 4294 5818 4350
rect 5886 4294 5942 4350
rect 5514 4170 5570 4226
rect 5638 4170 5694 4226
rect 5762 4170 5818 4226
rect 5886 4170 5942 4226
rect 5514 4046 5570 4102
rect 5638 4046 5694 4102
rect 5762 4046 5818 4102
rect 5886 4046 5942 4102
rect 5514 3922 5570 3978
rect 5638 3922 5694 3978
rect 5762 3922 5818 3978
rect 5886 3922 5942 3978
rect 5514 -216 5570 -160
rect 5638 -216 5694 -160
rect 5762 -216 5818 -160
rect 5886 -216 5942 -160
rect 5514 -340 5570 -284
rect 5638 -340 5694 -284
rect 5762 -340 5818 -284
rect 5886 -340 5942 -284
rect 5514 -464 5570 -408
rect 5638 -464 5694 -408
rect 5762 -464 5818 -408
rect 5886 -464 5942 -408
rect 5514 -588 5570 -532
rect 5638 -588 5694 -532
rect 5762 -588 5818 -532
rect 5886 -588 5942 -532
rect -1820 -1176 -1764 -1120
rect -1696 -1176 -1640 -1120
rect -1572 -1176 -1516 -1120
rect -1448 -1176 -1392 -1120
rect -1820 -1300 -1764 -1244
rect -1696 -1300 -1640 -1244
rect -1572 -1300 -1516 -1244
rect -1448 -1300 -1392 -1244
rect -1820 -1424 -1764 -1368
rect -1696 -1424 -1640 -1368
rect -1572 -1424 -1516 -1368
rect -1448 -1424 -1392 -1368
rect -1820 -1548 -1764 -1492
rect -1696 -1548 -1640 -1492
rect -1572 -1548 -1516 -1492
rect -1448 -1548 -1392 -1492
rect 36234 4294 36290 4350
rect 36358 4294 36414 4350
rect 36482 4294 36538 4350
rect 36606 4294 36662 4350
rect 36234 4170 36290 4226
rect 36358 4170 36414 4226
rect 36482 4170 36538 4226
rect 36606 4170 36662 4226
rect 36234 4046 36290 4102
rect 36358 4046 36414 4102
rect 36482 4046 36538 4102
rect 36606 4046 36662 4102
rect 36234 3922 36290 3978
rect 36358 3922 36414 3978
rect 36482 3922 36538 3978
rect 36606 3922 36662 3978
rect 36234 -216 36290 -160
rect 36358 -216 36414 -160
rect 36482 -216 36538 -160
rect 36606 -216 36662 -160
rect 36234 -340 36290 -284
rect 36358 -340 36414 -284
rect 36482 -340 36538 -284
rect 36606 -340 36662 -284
rect 36234 -464 36290 -408
rect 36358 -464 36414 -408
rect 36482 -464 36538 -408
rect 36606 -464 36662 -408
rect 36234 -588 36290 -532
rect 36358 -588 36414 -532
rect 36482 -588 36538 -532
rect 36606 -588 36662 -532
rect 66954 4294 67010 4350
rect 67078 4294 67134 4350
rect 67202 4294 67258 4350
rect 67326 4294 67382 4350
rect 66954 4170 67010 4226
rect 67078 4170 67134 4226
rect 67202 4170 67258 4226
rect 67326 4170 67382 4226
rect 66954 4046 67010 4102
rect 67078 4046 67134 4102
rect 67202 4046 67258 4102
rect 67326 4046 67382 4102
rect 66954 3922 67010 3978
rect 67078 3922 67134 3978
rect 67202 3922 67258 3978
rect 67326 3922 67382 3978
rect 66954 -216 67010 -160
rect 67078 -216 67134 -160
rect 67202 -216 67258 -160
rect 67326 -216 67382 -160
rect 66954 -340 67010 -284
rect 67078 -340 67134 -284
rect 67202 -340 67258 -284
rect 67326 -340 67382 -284
rect 66954 -464 67010 -408
rect 67078 -464 67134 -408
rect 67202 -464 67258 -408
rect 67326 -464 67382 -408
rect 66954 -588 67010 -532
rect 67078 -588 67134 -532
rect 67202 -588 67258 -532
rect 67326 -588 67382 -532
rect 97674 4294 97730 4350
rect 97798 4294 97854 4350
rect 97922 4294 97978 4350
rect 98046 4294 98102 4350
rect 97674 4170 97730 4226
rect 97798 4170 97854 4226
rect 97922 4170 97978 4226
rect 98046 4170 98102 4226
rect 97674 4046 97730 4102
rect 97798 4046 97854 4102
rect 97922 4046 97978 4102
rect 98046 4046 98102 4102
rect 97674 3922 97730 3978
rect 97798 3922 97854 3978
rect 97922 3922 97978 3978
rect 98046 3922 98102 3978
rect 97674 -216 97730 -160
rect 97798 -216 97854 -160
rect 97922 -216 97978 -160
rect 98046 -216 98102 -160
rect 97674 -340 97730 -284
rect 97798 -340 97854 -284
rect 97922 -340 97978 -284
rect 98046 -340 98102 -284
rect 97674 -464 97730 -408
rect 97798 -464 97854 -408
rect 97922 -464 97978 -408
rect 98046 -464 98102 -408
rect 97674 -588 97730 -532
rect 97798 -588 97854 -532
rect 97922 -588 97978 -532
rect 98046 -588 98102 -532
rect 128394 4294 128450 4350
rect 128518 4294 128574 4350
rect 128642 4294 128698 4350
rect 128766 4294 128822 4350
rect 128394 4170 128450 4226
rect 128518 4170 128574 4226
rect 128642 4170 128698 4226
rect 128766 4170 128822 4226
rect 128394 4046 128450 4102
rect 128518 4046 128574 4102
rect 128642 4046 128698 4102
rect 128766 4046 128822 4102
rect 128394 3922 128450 3978
rect 128518 3922 128574 3978
rect 128642 3922 128698 3978
rect 128766 3922 128822 3978
rect 128394 -216 128450 -160
rect 128518 -216 128574 -160
rect 128642 -216 128698 -160
rect 128766 -216 128822 -160
rect 128394 -340 128450 -284
rect 128518 -340 128574 -284
rect 128642 -340 128698 -284
rect 128766 -340 128822 -284
rect 128394 -464 128450 -408
rect 128518 -464 128574 -408
rect 128642 -464 128698 -408
rect 128766 -464 128822 -408
rect 128394 -588 128450 -532
rect 128518 -588 128574 -532
rect 128642 -588 128698 -532
rect 128766 -588 128822 -532
rect 159114 4294 159170 4350
rect 159238 4294 159294 4350
rect 159362 4294 159418 4350
rect 159486 4294 159542 4350
rect 159114 4170 159170 4226
rect 159238 4170 159294 4226
rect 159362 4170 159418 4226
rect 159486 4170 159542 4226
rect 159114 4046 159170 4102
rect 159238 4046 159294 4102
rect 159362 4046 159418 4102
rect 159486 4046 159542 4102
rect 159114 3922 159170 3978
rect 159238 3922 159294 3978
rect 159362 3922 159418 3978
rect 159486 3922 159542 3978
rect 159114 -216 159170 -160
rect 159238 -216 159294 -160
rect 159362 -216 159418 -160
rect 159486 -216 159542 -160
rect 159114 -340 159170 -284
rect 159238 -340 159294 -284
rect 159362 -340 159418 -284
rect 159486 -340 159542 -284
rect 159114 -464 159170 -408
rect 159238 -464 159294 -408
rect 159362 -464 159418 -408
rect 159486 -464 159542 -408
rect 159114 -588 159170 -532
rect 159238 -588 159294 -532
rect 159362 -588 159418 -532
rect 159486 -588 159542 -532
rect 189834 4294 189890 4350
rect 189958 4294 190014 4350
rect 190082 4294 190138 4350
rect 190206 4294 190262 4350
rect 189834 4170 189890 4226
rect 189958 4170 190014 4226
rect 190082 4170 190138 4226
rect 190206 4170 190262 4226
rect 189834 4046 189890 4102
rect 189958 4046 190014 4102
rect 190082 4046 190138 4102
rect 190206 4046 190262 4102
rect 189834 3922 189890 3978
rect 189958 3922 190014 3978
rect 190082 3922 190138 3978
rect 190206 3922 190262 3978
rect 189834 -216 189890 -160
rect 189958 -216 190014 -160
rect 190082 -216 190138 -160
rect 190206 -216 190262 -160
rect 189834 -340 189890 -284
rect 189958 -340 190014 -284
rect 190082 -340 190138 -284
rect 190206 -340 190262 -284
rect 189834 -464 189890 -408
rect 189958 -464 190014 -408
rect 190082 -464 190138 -408
rect 190206 -464 190262 -408
rect 189834 -588 189890 -532
rect 189958 -588 190014 -532
rect 190082 -588 190138 -532
rect 190206 -588 190262 -532
rect 220554 4294 220610 4350
rect 220678 4294 220734 4350
rect 220802 4294 220858 4350
rect 220926 4294 220982 4350
rect 220554 4170 220610 4226
rect 220678 4170 220734 4226
rect 220802 4170 220858 4226
rect 220926 4170 220982 4226
rect 220554 4046 220610 4102
rect 220678 4046 220734 4102
rect 220802 4046 220858 4102
rect 220926 4046 220982 4102
rect 220554 3922 220610 3978
rect 220678 3922 220734 3978
rect 220802 3922 220858 3978
rect 220926 3922 220982 3978
rect 220554 -216 220610 -160
rect 220678 -216 220734 -160
rect 220802 -216 220858 -160
rect 220926 -216 220982 -160
rect 220554 -340 220610 -284
rect 220678 -340 220734 -284
rect 220802 -340 220858 -284
rect 220926 -340 220982 -284
rect 220554 -464 220610 -408
rect 220678 -464 220734 -408
rect 220802 -464 220858 -408
rect 220926 -464 220982 -408
rect 220554 -588 220610 -532
rect 220678 -588 220734 -532
rect 220802 -588 220858 -532
rect 220926 -588 220982 -532
rect 251274 4294 251330 4350
rect 251398 4294 251454 4350
rect 251522 4294 251578 4350
rect 251646 4294 251702 4350
rect 251274 4170 251330 4226
rect 251398 4170 251454 4226
rect 251522 4170 251578 4226
rect 251646 4170 251702 4226
rect 251274 4046 251330 4102
rect 251398 4046 251454 4102
rect 251522 4046 251578 4102
rect 251646 4046 251702 4102
rect 251274 3922 251330 3978
rect 251398 3922 251454 3978
rect 251522 3922 251578 3978
rect 251646 3922 251702 3978
rect 251274 -216 251330 -160
rect 251398 -216 251454 -160
rect 251522 -216 251578 -160
rect 251646 -216 251702 -160
rect 251274 -340 251330 -284
rect 251398 -340 251454 -284
rect 251522 -340 251578 -284
rect 251646 -340 251702 -284
rect 251274 -464 251330 -408
rect 251398 -464 251454 -408
rect 251522 -464 251578 -408
rect 251646 -464 251702 -408
rect 251274 -588 251330 -532
rect 251398 -588 251454 -532
rect 251522 -588 251578 -532
rect 251646 -588 251702 -532
rect 281994 4294 282050 4350
rect 282118 4294 282174 4350
rect 282242 4294 282298 4350
rect 282366 4294 282422 4350
rect 281994 4170 282050 4226
rect 282118 4170 282174 4226
rect 282242 4170 282298 4226
rect 282366 4170 282422 4226
rect 281994 4046 282050 4102
rect 282118 4046 282174 4102
rect 282242 4046 282298 4102
rect 282366 4046 282422 4102
rect 281994 3922 282050 3978
rect 282118 3922 282174 3978
rect 282242 3922 282298 3978
rect 282366 3922 282422 3978
rect 281994 -216 282050 -160
rect 282118 -216 282174 -160
rect 282242 -216 282298 -160
rect 282366 -216 282422 -160
rect 281994 -340 282050 -284
rect 282118 -340 282174 -284
rect 282242 -340 282298 -284
rect 282366 -340 282422 -284
rect 281994 -464 282050 -408
rect 282118 -464 282174 -408
rect 282242 -464 282298 -408
rect 282366 -464 282422 -408
rect 281994 -588 282050 -532
rect 282118 -588 282174 -532
rect 282242 -588 282298 -532
rect 282366 -588 282422 -532
rect 312714 4294 312770 4350
rect 312838 4294 312894 4350
rect 312962 4294 313018 4350
rect 313086 4294 313142 4350
rect 312714 4170 312770 4226
rect 312838 4170 312894 4226
rect 312962 4170 313018 4226
rect 313086 4170 313142 4226
rect 312714 4046 312770 4102
rect 312838 4046 312894 4102
rect 312962 4046 313018 4102
rect 313086 4046 313142 4102
rect 312714 3922 312770 3978
rect 312838 3922 312894 3978
rect 312962 3922 313018 3978
rect 313086 3922 313142 3978
rect 312714 -216 312770 -160
rect 312838 -216 312894 -160
rect 312962 -216 313018 -160
rect 313086 -216 313142 -160
rect 312714 -340 312770 -284
rect 312838 -340 312894 -284
rect 312962 -340 313018 -284
rect 313086 -340 313142 -284
rect 312714 -464 312770 -408
rect 312838 -464 312894 -408
rect 312962 -464 313018 -408
rect 313086 -464 313142 -408
rect 312714 -588 312770 -532
rect 312838 -588 312894 -532
rect 312962 -588 313018 -532
rect 313086 -588 313142 -532
rect 343434 4294 343490 4350
rect 343558 4294 343614 4350
rect 343682 4294 343738 4350
rect 343806 4294 343862 4350
rect 343434 4170 343490 4226
rect 343558 4170 343614 4226
rect 343682 4170 343738 4226
rect 343806 4170 343862 4226
rect 343434 4046 343490 4102
rect 343558 4046 343614 4102
rect 343682 4046 343738 4102
rect 343806 4046 343862 4102
rect 343434 3922 343490 3978
rect 343558 3922 343614 3978
rect 343682 3922 343738 3978
rect 343806 3922 343862 3978
rect 343434 -216 343490 -160
rect 343558 -216 343614 -160
rect 343682 -216 343738 -160
rect 343806 -216 343862 -160
rect 343434 -340 343490 -284
rect 343558 -340 343614 -284
rect 343682 -340 343738 -284
rect 343806 -340 343862 -284
rect 343434 -464 343490 -408
rect 343558 -464 343614 -408
rect 343682 -464 343738 -408
rect 343806 -464 343862 -408
rect 343434 -588 343490 -532
rect 343558 -588 343614 -532
rect 343682 -588 343738 -532
rect 343806 -588 343862 -532
rect 374154 4294 374210 4350
rect 374278 4294 374334 4350
rect 374402 4294 374458 4350
rect 374526 4294 374582 4350
rect 374154 4170 374210 4226
rect 374278 4170 374334 4226
rect 374402 4170 374458 4226
rect 374526 4170 374582 4226
rect 374154 4046 374210 4102
rect 374278 4046 374334 4102
rect 374402 4046 374458 4102
rect 374526 4046 374582 4102
rect 374154 3922 374210 3978
rect 374278 3922 374334 3978
rect 374402 3922 374458 3978
rect 374526 3922 374582 3978
rect 374154 -216 374210 -160
rect 374278 -216 374334 -160
rect 374402 -216 374458 -160
rect 374526 -216 374582 -160
rect 374154 -340 374210 -284
rect 374278 -340 374334 -284
rect 374402 -340 374458 -284
rect 374526 -340 374582 -284
rect 374154 -464 374210 -408
rect 374278 -464 374334 -408
rect 374402 -464 374458 -408
rect 374526 -464 374582 -408
rect 374154 -588 374210 -532
rect 374278 -588 374334 -532
rect 374402 -588 374458 -532
rect 374526 -588 374582 -532
rect 404874 4294 404930 4350
rect 404998 4294 405054 4350
rect 405122 4294 405178 4350
rect 405246 4294 405302 4350
rect 404874 4170 404930 4226
rect 404998 4170 405054 4226
rect 405122 4170 405178 4226
rect 405246 4170 405302 4226
rect 404874 4046 404930 4102
rect 404998 4046 405054 4102
rect 405122 4046 405178 4102
rect 405246 4046 405302 4102
rect 404874 3922 404930 3978
rect 404998 3922 405054 3978
rect 405122 3922 405178 3978
rect 405246 3922 405302 3978
rect 404874 -216 404930 -160
rect 404998 -216 405054 -160
rect 405122 -216 405178 -160
rect 405246 -216 405302 -160
rect 404874 -340 404930 -284
rect 404998 -340 405054 -284
rect 405122 -340 405178 -284
rect 405246 -340 405302 -284
rect 404874 -464 404930 -408
rect 404998 -464 405054 -408
rect 405122 -464 405178 -408
rect 405246 -464 405302 -408
rect 404874 -588 404930 -532
rect 404998 -588 405054 -532
rect 405122 -588 405178 -532
rect 405246 -588 405302 -532
rect 435594 4294 435650 4350
rect 435718 4294 435774 4350
rect 435842 4294 435898 4350
rect 435966 4294 436022 4350
rect 435594 4170 435650 4226
rect 435718 4170 435774 4226
rect 435842 4170 435898 4226
rect 435966 4170 436022 4226
rect 435594 4046 435650 4102
rect 435718 4046 435774 4102
rect 435842 4046 435898 4102
rect 435966 4046 436022 4102
rect 435594 3922 435650 3978
rect 435718 3922 435774 3978
rect 435842 3922 435898 3978
rect 435966 3922 436022 3978
rect 435594 -216 435650 -160
rect 435718 -216 435774 -160
rect 435842 -216 435898 -160
rect 435966 -216 436022 -160
rect 435594 -340 435650 -284
rect 435718 -340 435774 -284
rect 435842 -340 435898 -284
rect 435966 -340 436022 -284
rect 435594 -464 435650 -408
rect 435718 -464 435774 -408
rect 435842 -464 435898 -408
rect 435966 -464 436022 -408
rect 435594 -588 435650 -532
rect 435718 -588 435774 -532
rect 435842 -588 435898 -532
rect 435966 -588 436022 -532
rect 466314 4294 466370 4350
rect 466438 4294 466494 4350
rect 466562 4294 466618 4350
rect 466686 4294 466742 4350
rect 466314 4170 466370 4226
rect 466438 4170 466494 4226
rect 466562 4170 466618 4226
rect 466686 4170 466742 4226
rect 466314 4046 466370 4102
rect 466438 4046 466494 4102
rect 466562 4046 466618 4102
rect 466686 4046 466742 4102
rect 466314 3922 466370 3978
rect 466438 3922 466494 3978
rect 466562 3922 466618 3978
rect 466686 3922 466742 3978
rect 466314 -216 466370 -160
rect 466438 -216 466494 -160
rect 466562 -216 466618 -160
rect 466686 -216 466742 -160
rect 466314 -340 466370 -284
rect 466438 -340 466494 -284
rect 466562 -340 466618 -284
rect 466686 -340 466742 -284
rect 466314 -464 466370 -408
rect 466438 -464 466494 -408
rect 466562 -464 466618 -408
rect 466686 -464 466742 -408
rect 466314 -588 466370 -532
rect 466438 -588 466494 -532
rect 466562 -588 466618 -532
rect 466686 -588 466742 -532
rect 497034 4294 497090 4350
rect 497158 4294 497214 4350
rect 497282 4294 497338 4350
rect 497406 4294 497462 4350
rect 497034 4170 497090 4226
rect 497158 4170 497214 4226
rect 497282 4170 497338 4226
rect 497406 4170 497462 4226
rect 497034 4046 497090 4102
rect 497158 4046 497214 4102
rect 497282 4046 497338 4102
rect 497406 4046 497462 4102
rect 497034 3922 497090 3978
rect 497158 3922 497214 3978
rect 497282 3922 497338 3978
rect 497406 3922 497462 3978
rect 497034 -216 497090 -160
rect 497158 -216 497214 -160
rect 497282 -216 497338 -160
rect 497406 -216 497462 -160
rect 497034 -340 497090 -284
rect 497158 -340 497214 -284
rect 497282 -340 497338 -284
rect 497406 -340 497462 -284
rect 497034 -464 497090 -408
rect 497158 -464 497214 -408
rect 497282 -464 497338 -408
rect 497406 -464 497462 -408
rect 497034 -588 497090 -532
rect 497158 -588 497214 -532
rect 497282 -588 497338 -532
rect 497406 -588 497462 -532
rect 557452 4922 557508 4978
rect 527754 4294 527810 4350
rect 527878 4294 527934 4350
rect 528002 4294 528058 4350
rect 528126 4294 528182 4350
rect 527754 4170 527810 4226
rect 527878 4170 527934 4226
rect 528002 4170 528058 4226
rect 528126 4170 528182 4226
rect 527754 4046 527810 4102
rect 527878 4046 527934 4102
rect 528002 4046 528058 4102
rect 528126 4046 528182 4102
rect 527754 3922 527810 3978
rect 527878 3922 527934 3978
rect 528002 3922 528058 3978
rect 528126 3922 528182 3978
rect 527754 -216 527810 -160
rect 527878 -216 527934 -160
rect 528002 -216 528058 -160
rect 528126 -216 528182 -160
rect 527754 -340 527810 -284
rect 527878 -340 527934 -284
rect 528002 -340 528058 -284
rect 528126 -340 528182 -284
rect 527754 -464 527810 -408
rect 527878 -464 527934 -408
rect 528002 -464 528058 -408
rect 528126 -464 528182 -408
rect 527754 -588 527810 -532
rect 527878 -588 527934 -532
rect 528002 -588 528058 -532
rect 528126 -588 528182 -532
rect 561036 4742 561092 4798
rect 576828 4922 576884 4978
rect 558474 4294 558530 4350
rect 558598 4294 558654 4350
rect 558722 4294 558778 4350
rect 558846 4294 558902 4350
rect 558474 4170 558530 4226
rect 558598 4170 558654 4226
rect 558722 4170 558778 4226
rect 558846 4170 558902 4226
rect 558474 4046 558530 4102
rect 558598 4046 558654 4102
rect 558722 4046 558778 4102
rect 558846 4046 558902 4102
rect 558474 3922 558530 3978
rect 558598 3922 558654 3978
rect 558722 3922 558778 3978
rect 558846 3922 558902 3978
rect 580636 4742 580692 4798
rect 589194 4294 589250 4350
rect 589318 4294 589374 4350
rect 589442 4294 589498 4350
rect 589566 4294 589622 4350
rect 589194 4170 589250 4226
rect 589318 4170 589374 4226
rect 589442 4170 589498 4226
rect 589566 4170 589622 4226
rect 589194 4046 589250 4102
rect 589318 4046 589374 4102
rect 589442 4046 589498 4102
rect 589566 4046 589622 4102
rect 589194 3922 589250 3978
rect 589318 3922 589374 3978
rect 589442 3922 589498 3978
rect 589566 3922 589622 3978
rect 558474 -216 558530 -160
rect 558598 -216 558654 -160
rect 558722 -216 558778 -160
rect 558846 -216 558902 -160
rect 558474 -340 558530 -284
rect 558598 -340 558654 -284
rect 558722 -340 558778 -284
rect 558846 -340 558902 -284
rect 558474 -464 558530 -408
rect 558598 -464 558654 -408
rect 558722 -464 558778 -408
rect 558846 -464 558902 -408
rect 558474 -588 558530 -532
rect 558598 -588 558654 -532
rect 558722 -588 558778 -532
rect 558846 -588 558902 -532
rect 589194 -216 589250 -160
rect 589318 -216 589374 -160
rect 589442 -216 589498 -160
rect 589566 -216 589622 -160
rect 589194 -340 589250 -284
rect 589318 -340 589374 -284
rect 589442 -340 589498 -284
rect 589566 -340 589622 -284
rect 589194 -464 589250 -408
rect 589318 -464 589374 -408
rect 589442 -464 589498 -408
rect 589566 -464 589622 -408
rect 589194 -588 589250 -532
rect 589318 -588 589374 -532
rect 589442 -588 589498 -532
rect 589566 -588 589622 -532
rect 592914 46294 592970 46350
rect 593038 46294 593094 46350
rect 593162 46294 593218 46350
rect 593286 46294 593342 46350
rect 592914 46170 592970 46226
rect 593038 46170 593094 46226
rect 593162 46170 593218 46226
rect 593286 46170 593342 46226
rect 592914 46046 592970 46102
rect 593038 46046 593094 46102
rect 593162 46046 593218 46102
rect 593286 46046 593342 46102
rect 592914 45922 592970 45978
rect 593038 45922 593094 45978
rect 593162 45922 593218 45978
rect 593286 45922 593342 45978
rect 592914 28294 592970 28350
rect 593038 28294 593094 28350
rect 593162 28294 593218 28350
rect 593286 28294 593342 28350
rect 592914 28170 592970 28226
rect 593038 28170 593094 28226
rect 593162 28170 593218 28226
rect 593286 28170 593342 28226
rect 592914 28046 592970 28102
rect 593038 28046 593094 28102
rect 593162 28046 593218 28102
rect 593286 28046 593342 28102
rect 592914 27922 592970 27978
rect 593038 27922 593094 27978
rect 593162 27922 593218 27978
rect 593286 27922 593342 27978
rect 592914 10294 592970 10350
rect 593038 10294 593094 10350
rect 593162 10294 593218 10350
rect 593286 10294 593342 10350
rect 592914 10170 592970 10226
rect 593038 10170 593094 10226
rect 593162 10170 593218 10226
rect 593286 10170 593342 10226
rect 592914 10046 592970 10102
rect 593038 10046 593094 10102
rect 593162 10046 593218 10102
rect 593286 10046 593342 10102
rect 592914 9922 592970 9978
rect 593038 9922 593094 9978
rect 593162 9922 593218 9978
rect 593286 9922 593342 9978
rect 596496 597156 596552 597212
rect 596620 597156 596676 597212
rect 596744 597156 596800 597212
rect 596868 597156 596924 597212
rect 596496 597032 596552 597088
rect 596620 597032 596676 597088
rect 596744 597032 596800 597088
rect 596868 597032 596924 597088
rect 596496 596908 596552 596964
rect 596620 596908 596676 596964
rect 596744 596908 596800 596964
rect 596868 596908 596924 596964
rect 596496 596784 596552 596840
rect 596620 596784 596676 596840
rect 596744 596784 596800 596840
rect 596868 596784 596924 596840
rect 596496 580294 596552 580350
rect 596620 580294 596676 580350
rect 596744 580294 596800 580350
rect 596868 580294 596924 580350
rect 596496 580170 596552 580226
rect 596620 580170 596676 580226
rect 596744 580170 596800 580226
rect 596868 580170 596924 580226
rect 596496 580046 596552 580102
rect 596620 580046 596676 580102
rect 596744 580046 596800 580102
rect 596868 580046 596924 580102
rect 596496 579922 596552 579978
rect 596620 579922 596676 579978
rect 596744 579922 596800 579978
rect 596868 579922 596924 579978
rect 596496 562294 596552 562350
rect 596620 562294 596676 562350
rect 596744 562294 596800 562350
rect 596868 562294 596924 562350
rect 596496 562170 596552 562226
rect 596620 562170 596676 562226
rect 596744 562170 596800 562226
rect 596868 562170 596924 562226
rect 596496 562046 596552 562102
rect 596620 562046 596676 562102
rect 596744 562046 596800 562102
rect 596868 562046 596924 562102
rect 596496 561922 596552 561978
rect 596620 561922 596676 561978
rect 596744 561922 596800 561978
rect 596868 561922 596924 561978
rect 596496 544294 596552 544350
rect 596620 544294 596676 544350
rect 596744 544294 596800 544350
rect 596868 544294 596924 544350
rect 596496 544170 596552 544226
rect 596620 544170 596676 544226
rect 596744 544170 596800 544226
rect 596868 544170 596924 544226
rect 596496 544046 596552 544102
rect 596620 544046 596676 544102
rect 596744 544046 596800 544102
rect 596868 544046 596924 544102
rect 596496 543922 596552 543978
rect 596620 543922 596676 543978
rect 596744 543922 596800 543978
rect 596868 543922 596924 543978
rect 596496 526294 596552 526350
rect 596620 526294 596676 526350
rect 596744 526294 596800 526350
rect 596868 526294 596924 526350
rect 596496 526170 596552 526226
rect 596620 526170 596676 526226
rect 596744 526170 596800 526226
rect 596868 526170 596924 526226
rect 596496 526046 596552 526102
rect 596620 526046 596676 526102
rect 596744 526046 596800 526102
rect 596868 526046 596924 526102
rect 596496 525922 596552 525978
rect 596620 525922 596676 525978
rect 596744 525922 596800 525978
rect 596868 525922 596924 525978
rect 596496 508294 596552 508350
rect 596620 508294 596676 508350
rect 596744 508294 596800 508350
rect 596868 508294 596924 508350
rect 596496 508170 596552 508226
rect 596620 508170 596676 508226
rect 596744 508170 596800 508226
rect 596868 508170 596924 508226
rect 596496 508046 596552 508102
rect 596620 508046 596676 508102
rect 596744 508046 596800 508102
rect 596868 508046 596924 508102
rect 596496 507922 596552 507978
rect 596620 507922 596676 507978
rect 596744 507922 596800 507978
rect 596868 507922 596924 507978
rect 596496 490294 596552 490350
rect 596620 490294 596676 490350
rect 596744 490294 596800 490350
rect 596868 490294 596924 490350
rect 596496 490170 596552 490226
rect 596620 490170 596676 490226
rect 596744 490170 596800 490226
rect 596868 490170 596924 490226
rect 596496 490046 596552 490102
rect 596620 490046 596676 490102
rect 596744 490046 596800 490102
rect 596868 490046 596924 490102
rect 596496 489922 596552 489978
rect 596620 489922 596676 489978
rect 596744 489922 596800 489978
rect 596868 489922 596924 489978
rect 596496 472294 596552 472350
rect 596620 472294 596676 472350
rect 596744 472294 596800 472350
rect 596868 472294 596924 472350
rect 596496 472170 596552 472226
rect 596620 472170 596676 472226
rect 596744 472170 596800 472226
rect 596868 472170 596924 472226
rect 596496 472046 596552 472102
rect 596620 472046 596676 472102
rect 596744 472046 596800 472102
rect 596868 472046 596924 472102
rect 596496 471922 596552 471978
rect 596620 471922 596676 471978
rect 596744 471922 596800 471978
rect 596868 471922 596924 471978
rect 596496 454294 596552 454350
rect 596620 454294 596676 454350
rect 596744 454294 596800 454350
rect 596868 454294 596924 454350
rect 596496 454170 596552 454226
rect 596620 454170 596676 454226
rect 596744 454170 596800 454226
rect 596868 454170 596924 454226
rect 596496 454046 596552 454102
rect 596620 454046 596676 454102
rect 596744 454046 596800 454102
rect 596868 454046 596924 454102
rect 596496 453922 596552 453978
rect 596620 453922 596676 453978
rect 596744 453922 596800 453978
rect 596868 453922 596924 453978
rect 596496 436294 596552 436350
rect 596620 436294 596676 436350
rect 596744 436294 596800 436350
rect 596868 436294 596924 436350
rect 596496 436170 596552 436226
rect 596620 436170 596676 436226
rect 596744 436170 596800 436226
rect 596868 436170 596924 436226
rect 596496 436046 596552 436102
rect 596620 436046 596676 436102
rect 596744 436046 596800 436102
rect 596868 436046 596924 436102
rect 596496 435922 596552 435978
rect 596620 435922 596676 435978
rect 596744 435922 596800 435978
rect 596868 435922 596924 435978
rect 596496 418294 596552 418350
rect 596620 418294 596676 418350
rect 596744 418294 596800 418350
rect 596868 418294 596924 418350
rect 596496 418170 596552 418226
rect 596620 418170 596676 418226
rect 596744 418170 596800 418226
rect 596868 418170 596924 418226
rect 596496 418046 596552 418102
rect 596620 418046 596676 418102
rect 596744 418046 596800 418102
rect 596868 418046 596924 418102
rect 596496 417922 596552 417978
rect 596620 417922 596676 417978
rect 596744 417922 596800 417978
rect 596868 417922 596924 417978
rect 596496 400294 596552 400350
rect 596620 400294 596676 400350
rect 596744 400294 596800 400350
rect 596868 400294 596924 400350
rect 596496 400170 596552 400226
rect 596620 400170 596676 400226
rect 596744 400170 596800 400226
rect 596868 400170 596924 400226
rect 596496 400046 596552 400102
rect 596620 400046 596676 400102
rect 596744 400046 596800 400102
rect 596868 400046 596924 400102
rect 596496 399922 596552 399978
rect 596620 399922 596676 399978
rect 596744 399922 596800 399978
rect 596868 399922 596924 399978
rect 596496 382294 596552 382350
rect 596620 382294 596676 382350
rect 596744 382294 596800 382350
rect 596868 382294 596924 382350
rect 596496 382170 596552 382226
rect 596620 382170 596676 382226
rect 596744 382170 596800 382226
rect 596868 382170 596924 382226
rect 596496 382046 596552 382102
rect 596620 382046 596676 382102
rect 596744 382046 596800 382102
rect 596868 382046 596924 382102
rect 596496 381922 596552 381978
rect 596620 381922 596676 381978
rect 596744 381922 596800 381978
rect 596868 381922 596924 381978
rect 596496 364294 596552 364350
rect 596620 364294 596676 364350
rect 596744 364294 596800 364350
rect 596868 364294 596924 364350
rect 596496 364170 596552 364226
rect 596620 364170 596676 364226
rect 596744 364170 596800 364226
rect 596868 364170 596924 364226
rect 596496 364046 596552 364102
rect 596620 364046 596676 364102
rect 596744 364046 596800 364102
rect 596868 364046 596924 364102
rect 596496 363922 596552 363978
rect 596620 363922 596676 363978
rect 596744 363922 596800 363978
rect 596868 363922 596924 363978
rect 596496 346294 596552 346350
rect 596620 346294 596676 346350
rect 596744 346294 596800 346350
rect 596868 346294 596924 346350
rect 596496 346170 596552 346226
rect 596620 346170 596676 346226
rect 596744 346170 596800 346226
rect 596868 346170 596924 346226
rect 596496 346046 596552 346102
rect 596620 346046 596676 346102
rect 596744 346046 596800 346102
rect 596868 346046 596924 346102
rect 596496 345922 596552 345978
rect 596620 345922 596676 345978
rect 596744 345922 596800 345978
rect 596868 345922 596924 345978
rect 596496 328294 596552 328350
rect 596620 328294 596676 328350
rect 596744 328294 596800 328350
rect 596868 328294 596924 328350
rect 596496 328170 596552 328226
rect 596620 328170 596676 328226
rect 596744 328170 596800 328226
rect 596868 328170 596924 328226
rect 596496 328046 596552 328102
rect 596620 328046 596676 328102
rect 596744 328046 596800 328102
rect 596868 328046 596924 328102
rect 596496 327922 596552 327978
rect 596620 327922 596676 327978
rect 596744 327922 596800 327978
rect 596868 327922 596924 327978
rect 596496 310294 596552 310350
rect 596620 310294 596676 310350
rect 596744 310294 596800 310350
rect 596868 310294 596924 310350
rect 596496 310170 596552 310226
rect 596620 310170 596676 310226
rect 596744 310170 596800 310226
rect 596868 310170 596924 310226
rect 596496 310046 596552 310102
rect 596620 310046 596676 310102
rect 596744 310046 596800 310102
rect 596868 310046 596924 310102
rect 596496 309922 596552 309978
rect 596620 309922 596676 309978
rect 596744 309922 596800 309978
rect 596868 309922 596924 309978
rect 596496 292294 596552 292350
rect 596620 292294 596676 292350
rect 596744 292294 596800 292350
rect 596868 292294 596924 292350
rect 596496 292170 596552 292226
rect 596620 292170 596676 292226
rect 596744 292170 596800 292226
rect 596868 292170 596924 292226
rect 596496 292046 596552 292102
rect 596620 292046 596676 292102
rect 596744 292046 596800 292102
rect 596868 292046 596924 292102
rect 596496 291922 596552 291978
rect 596620 291922 596676 291978
rect 596744 291922 596800 291978
rect 596868 291922 596924 291978
rect 596496 274294 596552 274350
rect 596620 274294 596676 274350
rect 596744 274294 596800 274350
rect 596868 274294 596924 274350
rect 596496 274170 596552 274226
rect 596620 274170 596676 274226
rect 596744 274170 596800 274226
rect 596868 274170 596924 274226
rect 596496 274046 596552 274102
rect 596620 274046 596676 274102
rect 596744 274046 596800 274102
rect 596868 274046 596924 274102
rect 596496 273922 596552 273978
rect 596620 273922 596676 273978
rect 596744 273922 596800 273978
rect 596868 273922 596924 273978
rect 596496 256294 596552 256350
rect 596620 256294 596676 256350
rect 596744 256294 596800 256350
rect 596868 256294 596924 256350
rect 596496 256170 596552 256226
rect 596620 256170 596676 256226
rect 596744 256170 596800 256226
rect 596868 256170 596924 256226
rect 596496 256046 596552 256102
rect 596620 256046 596676 256102
rect 596744 256046 596800 256102
rect 596868 256046 596924 256102
rect 596496 255922 596552 255978
rect 596620 255922 596676 255978
rect 596744 255922 596800 255978
rect 596868 255922 596924 255978
rect 596496 238294 596552 238350
rect 596620 238294 596676 238350
rect 596744 238294 596800 238350
rect 596868 238294 596924 238350
rect 596496 238170 596552 238226
rect 596620 238170 596676 238226
rect 596744 238170 596800 238226
rect 596868 238170 596924 238226
rect 596496 238046 596552 238102
rect 596620 238046 596676 238102
rect 596744 238046 596800 238102
rect 596868 238046 596924 238102
rect 596496 237922 596552 237978
rect 596620 237922 596676 237978
rect 596744 237922 596800 237978
rect 596868 237922 596924 237978
rect 596496 220294 596552 220350
rect 596620 220294 596676 220350
rect 596744 220294 596800 220350
rect 596868 220294 596924 220350
rect 596496 220170 596552 220226
rect 596620 220170 596676 220226
rect 596744 220170 596800 220226
rect 596868 220170 596924 220226
rect 596496 220046 596552 220102
rect 596620 220046 596676 220102
rect 596744 220046 596800 220102
rect 596868 220046 596924 220102
rect 596496 219922 596552 219978
rect 596620 219922 596676 219978
rect 596744 219922 596800 219978
rect 596868 219922 596924 219978
rect 596496 202294 596552 202350
rect 596620 202294 596676 202350
rect 596744 202294 596800 202350
rect 596868 202294 596924 202350
rect 596496 202170 596552 202226
rect 596620 202170 596676 202226
rect 596744 202170 596800 202226
rect 596868 202170 596924 202226
rect 596496 202046 596552 202102
rect 596620 202046 596676 202102
rect 596744 202046 596800 202102
rect 596868 202046 596924 202102
rect 596496 201922 596552 201978
rect 596620 201922 596676 201978
rect 596744 201922 596800 201978
rect 596868 201922 596924 201978
rect 596496 184294 596552 184350
rect 596620 184294 596676 184350
rect 596744 184294 596800 184350
rect 596868 184294 596924 184350
rect 596496 184170 596552 184226
rect 596620 184170 596676 184226
rect 596744 184170 596800 184226
rect 596868 184170 596924 184226
rect 596496 184046 596552 184102
rect 596620 184046 596676 184102
rect 596744 184046 596800 184102
rect 596868 184046 596924 184102
rect 596496 183922 596552 183978
rect 596620 183922 596676 183978
rect 596744 183922 596800 183978
rect 596868 183922 596924 183978
rect 596496 166294 596552 166350
rect 596620 166294 596676 166350
rect 596744 166294 596800 166350
rect 596868 166294 596924 166350
rect 596496 166170 596552 166226
rect 596620 166170 596676 166226
rect 596744 166170 596800 166226
rect 596868 166170 596924 166226
rect 596496 166046 596552 166102
rect 596620 166046 596676 166102
rect 596744 166046 596800 166102
rect 596868 166046 596924 166102
rect 596496 165922 596552 165978
rect 596620 165922 596676 165978
rect 596744 165922 596800 165978
rect 596868 165922 596924 165978
rect 596496 148294 596552 148350
rect 596620 148294 596676 148350
rect 596744 148294 596800 148350
rect 596868 148294 596924 148350
rect 596496 148170 596552 148226
rect 596620 148170 596676 148226
rect 596744 148170 596800 148226
rect 596868 148170 596924 148226
rect 596496 148046 596552 148102
rect 596620 148046 596676 148102
rect 596744 148046 596800 148102
rect 596868 148046 596924 148102
rect 596496 147922 596552 147978
rect 596620 147922 596676 147978
rect 596744 147922 596800 147978
rect 596868 147922 596924 147978
rect 596496 130294 596552 130350
rect 596620 130294 596676 130350
rect 596744 130294 596800 130350
rect 596868 130294 596924 130350
rect 596496 130170 596552 130226
rect 596620 130170 596676 130226
rect 596744 130170 596800 130226
rect 596868 130170 596924 130226
rect 596496 130046 596552 130102
rect 596620 130046 596676 130102
rect 596744 130046 596800 130102
rect 596868 130046 596924 130102
rect 596496 129922 596552 129978
rect 596620 129922 596676 129978
rect 596744 129922 596800 129978
rect 596868 129922 596924 129978
rect 596496 112294 596552 112350
rect 596620 112294 596676 112350
rect 596744 112294 596800 112350
rect 596868 112294 596924 112350
rect 596496 112170 596552 112226
rect 596620 112170 596676 112226
rect 596744 112170 596800 112226
rect 596868 112170 596924 112226
rect 596496 112046 596552 112102
rect 596620 112046 596676 112102
rect 596744 112046 596800 112102
rect 596868 112046 596924 112102
rect 596496 111922 596552 111978
rect 596620 111922 596676 111978
rect 596744 111922 596800 111978
rect 596868 111922 596924 111978
rect 596496 94294 596552 94350
rect 596620 94294 596676 94350
rect 596744 94294 596800 94350
rect 596868 94294 596924 94350
rect 596496 94170 596552 94226
rect 596620 94170 596676 94226
rect 596744 94170 596800 94226
rect 596868 94170 596924 94226
rect 596496 94046 596552 94102
rect 596620 94046 596676 94102
rect 596744 94046 596800 94102
rect 596868 94046 596924 94102
rect 596496 93922 596552 93978
rect 596620 93922 596676 93978
rect 596744 93922 596800 93978
rect 596868 93922 596924 93978
rect 596496 76294 596552 76350
rect 596620 76294 596676 76350
rect 596744 76294 596800 76350
rect 596868 76294 596924 76350
rect 596496 76170 596552 76226
rect 596620 76170 596676 76226
rect 596744 76170 596800 76226
rect 596868 76170 596924 76226
rect 596496 76046 596552 76102
rect 596620 76046 596676 76102
rect 596744 76046 596800 76102
rect 596868 76046 596924 76102
rect 596496 75922 596552 75978
rect 596620 75922 596676 75978
rect 596744 75922 596800 75978
rect 596868 75922 596924 75978
rect 596496 58294 596552 58350
rect 596620 58294 596676 58350
rect 596744 58294 596800 58350
rect 596868 58294 596924 58350
rect 596496 58170 596552 58226
rect 596620 58170 596676 58226
rect 596744 58170 596800 58226
rect 596868 58170 596924 58226
rect 596496 58046 596552 58102
rect 596620 58046 596676 58102
rect 596744 58046 596800 58102
rect 596868 58046 596924 58102
rect 596496 57922 596552 57978
rect 596620 57922 596676 57978
rect 596744 57922 596800 57978
rect 596868 57922 596924 57978
rect 596496 40294 596552 40350
rect 596620 40294 596676 40350
rect 596744 40294 596800 40350
rect 596868 40294 596924 40350
rect 596496 40170 596552 40226
rect 596620 40170 596676 40226
rect 596744 40170 596800 40226
rect 596868 40170 596924 40226
rect 596496 40046 596552 40102
rect 596620 40046 596676 40102
rect 596744 40046 596800 40102
rect 596868 40046 596924 40102
rect 596496 39922 596552 39978
rect 596620 39922 596676 39978
rect 596744 39922 596800 39978
rect 596868 39922 596924 39978
rect 596496 22294 596552 22350
rect 596620 22294 596676 22350
rect 596744 22294 596800 22350
rect 596868 22294 596924 22350
rect 596496 22170 596552 22226
rect 596620 22170 596676 22226
rect 596744 22170 596800 22226
rect 596868 22170 596924 22226
rect 596496 22046 596552 22102
rect 596620 22046 596676 22102
rect 596744 22046 596800 22102
rect 596868 22046 596924 22102
rect 596496 21922 596552 21978
rect 596620 21922 596676 21978
rect 596744 21922 596800 21978
rect 596868 21922 596924 21978
rect 596496 4294 596552 4350
rect 596620 4294 596676 4350
rect 596744 4294 596800 4350
rect 596868 4294 596924 4350
rect 596496 4170 596552 4226
rect 596620 4170 596676 4226
rect 596744 4170 596800 4226
rect 596868 4170 596924 4226
rect 596496 4046 596552 4102
rect 596620 4046 596676 4102
rect 596744 4046 596800 4102
rect 596868 4046 596924 4102
rect 596496 3922 596552 3978
rect 596620 3922 596676 3978
rect 596744 3922 596800 3978
rect 596868 3922 596924 3978
rect 596496 -216 596552 -160
rect 596620 -216 596676 -160
rect 596744 -216 596800 -160
rect 596868 -216 596924 -160
rect 596496 -340 596552 -284
rect 596620 -340 596676 -284
rect 596744 -340 596800 -284
rect 596868 -340 596924 -284
rect 596496 -464 596552 -408
rect 596620 -464 596676 -408
rect 596744 -464 596800 -408
rect 596868 -464 596924 -408
rect 596496 -588 596552 -532
rect 596620 -588 596676 -532
rect 596744 -588 596800 -532
rect 596868 -588 596924 -532
rect 597456 586294 597512 586350
rect 597580 586294 597636 586350
rect 597704 586294 597760 586350
rect 597828 586294 597884 586350
rect 597456 586170 597512 586226
rect 597580 586170 597636 586226
rect 597704 586170 597760 586226
rect 597828 586170 597884 586226
rect 597456 586046 597512 586102
rect 597580 586046 597636 586102
rect 597704 586046 597760 586102
rect 597828 586046 597884 586102
rect 597456 585922 597512 585978
rect 597580 585922 597636 585978
rect 597704 585922 597760 585978
rect 597828 585922 597884 585978
rect 597456 568294 597512 568350
rect 597580 568294 597636 568350
rect 597704 568294 597760 568350
rect 597828 568294 597884 568350
rect 597456 568170 597512 568226
rect 597580 568170 597636 568226
rect 597704 568170 597760 568226
rect 597828 568170 597884 568226
rect 597456 568046 597512 568102
rect 597580 568046 597636 568102
rect 597704 568046 597760 568102
rect 597828 568046 597884 568102
rect 597456 567922 597512 567978
rect 597580 567922 597636 567978
rect 597704 567922 597760 567978
rect 597828 567922 597884 567978
rect 597456 550294 597512 550350
rect 597580 550294 597636 550350
rect 597704 550294 597760 550350
rect 597828 550294 597884 550350
rect 597456 550170 597512 550226
rect 597580 550170 597636 550226
rect 597704 550170 597760 550226
rect 597828 550170 597884 550226
rect 597456 550046 597512 550102
rect 597580 550046 597636 550102
rect 597704 550046 597760 550102
rect 597828 550046 597884 550102
rect 597456 549922 597512 549978
rect 597580 549922 597636 549978
rect 597704 549922 597760 549978
rect 597828 549922 597884 549978
rect 597456 532294 597512 532350
rect 597580 532294 597636 532350
rect 597704 532294 597760 532350
rect 597828 532294 597884 532350
rect 597456 532170 597512 532226
rect 597580 532170 597636 532226
rect 597704 532170 597760 532226
rect 597828 532170 597884 532226
rect 597456 532046 597512 532102
rect 597580 532046 597636 532102
rect 597704 532046 597760 532102
rect 597828 532046 597884 532102
rect 597456 531922 597512 531978
rect 597580 531922 597636 531978
rect 597704 531922 597760 531978
rect 597828 531922 597884 531978
rect 597456 514294 597512 514350
rect 597580 514294 597636 514350
rect 597704 514294 597760 514350
rect 597828 514294 597884 514350
rect 597456 514170 597512 514226
rect 597580 514170 597636 514226
rect 597704 514170 597760 514226
rect 597828 514170 597884 514226
rect 597456 514046 597512 514102
rect 597580 514046 597636 514102
rect 597704 514046 597760 514102
rect 597828 514046 597884 514102
rect 597456 513922 597512 513978
rect 597580 513922 597636 513978
rect 597704 513922 597760 513978
rect 597828 513922 597884 513978
rect 597456 496294 597512 496350
rect 597580 496294 597636 496350
rect 597704 496294 597760 496350
rect 597828 496294 597884 496350
rect 597456 496170 597512 496226
rect 597580 496170 597636 496226
rect 597704 496170 597760 496226
rect 597828 496170 597884 496226
rect 597456 496046 597512 496102
rect 597580 496046 597636 496102
rect 597704 496046 597760 496102
rect 597828 496046 597884 496102
rect 597456 495922 597512 495978
rect 597580 495922 597636 495978
rect 597704 495922 597760 495978
rect 597828 495922 597884 495978
rect 597456 478294 597512 478350
rect 597580 478294 597636 478350
rect 597704 478294 597760 478350
rect 597828 478294 597884 478350
rect 597456 478170 597512 478226
rect 597580 478170 597636 478226
rect 597704 478170 597760 478226
rect 597828 478170 597884 478226
rect 597456 478046 597512 478102
rect 597580 478046 597636 478102
rect 597704 478046 597760 478102
rect 597828 478046 597884 478102
rect 597456 477922 597512 477978
rect 597580 477922 597636 477978
rect 597704 477922 597760 477978
rect 597828 477922 597884 477978
rect 597456 460294 597512 460350
rect 597580 460294 597636 460350
rect 597704 460294 597760 460350
rect 597828 460294 597884 460350
rect 597456 460170 597512 460226
rect 597580 460170 597636 460226
rect 597704 460170 597760 460226
rect 597828 460170 597884 460226
rect 597456 460046 597512 460102
rect 597580 460046 597636 460102
rect 597704 460046 597760 460102
rect 597828 460046 597884 460102
rect 597456 459922 597512 459978
rect 597580 459922 597636 459978
rect 597704 459922 597760 459978
rect 597828 459922 597884 459978
rect 597456 442294 597512 442350
rect 597580 442294 597636 442350
rect 597704 442294 597760 442350
rect 597828 442294 597884 442350
rect 597456 442170 597512 442226
rect 597580 442170 597636 442226
rect 597704 442170 597760 442226
rect 597828 442170 597884 442226
rect 597456 442046 597512 442102
rect 597580 442046 597636 442102
rect 597704 442046 597760 442102
rect 597828 442046 597884 442102
rect 597456 441922 597512 441978
rect 597580 441922 597636 441978
rect 597704 441922 597760 441978
rect 597828 441922 597884 441978
rect 597456 424294 597512 424350
rect 597580 424294 597636 424350
rect 597704 424294 597760 424350
rect 597828 424294 597884 424350
rect 597456 424170 597512 424226
rect 597580 424170 597636 424226
rect 597704 424170 597760 424226
rect 597828 424170 597884 424226
rect 597456 424046 597512 424102
rect 597580 424046 597636 424102
rect 597704 424046 597760 424102
rect 597828 424046 597884 424102
rect 597456 423922 597512 423978
rect 597580 423922 597636 423978
rect 597704 423922 597760 423978
rect 597828 423922 597884 423978
rect 597456 406294 597512 406350
rect 597580 406294 597636 406350
rect 597704 406294 597760 406350
rect 597828 406294 597884 406350
rect 597456 406170 597512 406226
rect 597580 406170 597636 406226
rect 597704 406170 597760 406226
rect 597828 406170 597884 406226
rect 597456 406046 597512 406102
rect 597580 406046 597636 406102
rect 597704 406046 597760 406102
rect 597828 406046 597884 406102
rect 597456 405922 597512 405978
rect 597580 405922 597636 405978
rect 597704 405922 597760 405978
rect 597828 405922 597884 405978
rect 597456 388294 597512 388350
rect 597580 388294 597636 388350
rect 597704 388294 597760 388350
rect 597828 388294 597884 388350
rect 597456 388170 597512 388226
rect 597580 388170 597636 388226
rect 597704 388170 597760 388226
rect 597828 388170 597884 388226
rect 597456 388046 597512 388102
rect 597580 388046 597636 388102
rect 597704 388046 597760 388102
rect 597828 388046 597884 388102
rect 597456 387922 597512 387978
rect 597580 387922 597636 387978
rect 597704 387922 597760 387978
rect 597828 387922 597884 387978
rect 597456 370294 597512 370350
rect 597580 370294 597636 370350
rect 597704 370294 597760 370350
rect 597828 370294 597884 370350
rect 597456 370170 597512 370226
rect 597580 370170 597636 370226
rect 597704 370170 597760 370226
rect 597828 370170 597884 370226
rect 597456 370046 597512 370102
rect 597580 370046 597636 370102
rect 597704 370046 597760 370102
rect 597828 370046 597884 370102
rect 597456 369922 597512 369978
rect 597580 369922 597636 369978
rect 597704 369922 597760 369978
rect 597828 369922 597884 369978
rect 597456 352294 597512 352350
rect 597580 352294 597636 352350
rect 597704 352294 597760 352350
rect 597828 352294 597884 352350
rect 597456 352170 597512 352226
rect 597580 352170 597636 352226
rect 597704 352170 597760 352226
rect 597828 352170 597884 352226
rect 597456 352046 597512 352102
rect 597580 352046 597636 352102
rect 597704 352046 597760 352102
rect 597828 352046 597884 352102
rect 597456 351922 597512 351978
rect 597580 351922 597636 351978
rect 597704 351922 597760 351978
rect 597828 351922 597884 351978
rect 597456 334294 597512 334350
rect 597580 334294 597636 334350
rect 597704 334294 597760 334350
rect 597828 334294 597884 334350
rect 597456 334170 597512 334226
rect 597580 334170 597636 334226
rect 597704 334170 597760 334226
rect 597828 334170 597884 334226
rect 597456 334046 597512 334102
rect 597580 334046 597636 334102
rect 597704 334046 597760 334102
rect 597828 334046 597884 334102
rect 597456 333922 597512 333978
rect 597580 333922 597636 333978
rect 597704 333922 597760 333978
rect 597828 333922 597884 333978
rect 597456 316294 597512 316350
rect 597580 316294 597636 316350
rect 597704 316294 597760 316350
rect 597828 316294 597884 316350
rect 597456 316170 597512 316226
rect 597580 316170 597636 316226
rect 597704 316170 597760 316226
rect 597828 316170 597884 316226
rect 597456 316046 597512 316102
rect 597580 316046 597636 316102
rect 597704 316046 597760 316102
rect 597828 316046 597884 316102
rect 597456 315922 597512 315978
rect 597580 315922 597636 315978
rect 597704 315922 597760 315978
rect 597828 315922 597884 315978
rect 597456 298294 597512 298350
rect 597580 298294 597636 298350
rect 597704 298294 597760 298350
rect 597828 298294 597884 298350
rect 597456 298170 597512 298226
rect 597580 298170 597636 298226
rect 597704 298170 597760 298226
rect 597828 298170 597884 298226
rect 597456 298046 597512 298102
rect 597580 298046 597636 298102
rect 597704 298046 597760 298102
rect 597828 298046 597884 298102
rect 597456 297922 597512 297978
rect 597580 297922 597636 297978
rect 597704 297922 597760 297978
rect 597828 297922 597884 297978
rect 597456 280294 597512 280350
rect 597580 280294 597636 280350
rect 597704 280294 597760 280350
rect 597828 280294 597884 280350
rect 597456 280170 597512 280226
rect 597580 280170 597636 280226
rect 597704 280170 597760 280226
rect 597828 280170 597884 280226
rect 597456 280046 597512 280102
rect 597580 280046 597636 280102
rect 597704 280046 597760 280102
rect 597828 280046 597884 280102
rect 597456 279922 597512 279978
rect 597580 279922 597636 279978
rect 597704 279922 597760 279978
rect 597828 279922 597884 279978
rect 597456 262294 597512 262350
rect 597580 262294 597636 262350
rect 597704 262294 597760 262350
rect 597828 262294 597884 262350
rect 597456 262170 597512 262226
rect 597580 262170 597636 262226
rect 597704 262170 597760 262226
rect 597828 262170 597884 262226
rect 597456 262046 597512 262102
rect 597580 262046 597636 262102
rect 597704 262046 597760 262102
rect 597828 262046 597884 262102
rect 597456 261922 597512 261978
rect 597580 261922 597636 261978
rect 597704 261922 597760 261978
rect 597828 261922 597884 261978
rect 597456 244294 597512 244350
rect 597580 244294 597636 244350
rect 597704 244294 597760 244350
rect 597828 244294 597884 244350
rect 597456 244170 597512 244226
rect 597580 244170 597636 244226
rect 597704 244170 597760 244226
rect 597828 244170 597884 244226
rect 597456 244046 597512 244102
rect 597580 244046 597636 244102
rect 597704 244046 597760 244102
rect 597828 244046 597884 244102
rect 597456 243922 597512 243978
rect 597580 243922 597636 243978
rect 597704 243922 597760 243978
rect 597828 243922 597884 243978
rect 597456 226294 597512 226350
rect 597580 226294 597636 226350
rect 597704 226294 597760 226350
rect 597828 226294 597884 226350
rect 597456 226170 597512 226226
rect 597580 226170 597636 226226
rect 597704 226170 597760 226226
rect 597828 226170 597884 226226
rect 597456 226046 597512 226102
rect 597580 226046 597636 226102
rect 597704 226046 597760 226102
rect 597828 226046 597884 226102
rect 597456 225922 597512 225978
rect 597580 225922 597636 225978
rect 597704 225922 597760 225978
rect 597828 225922 597884 225978
rect 597456 208294 597512 208350
rect 597580 208294 597636 208350
rect 597704 208294 597760 208350
rect 597828 208294 597884 208350
rect 597456 208170 597512 208226
rect 597580 208170 597636 208226
rect 597704 208170 597760 208226
rect 597828 208170 597884 208226
rect 597456 208046 597512 208102
rect 597580 208046 597636 208102
rect 597704 208046 597760 208102
rect 597828 208046 597884 208102
rect 597456 207922 597512 207978
rect 597580 207922 597636 207978
rect 597704 207922 597760 207978
rect 597828 207922 597884 207978
rect 597456 190294 597512 190350
rect 597580 190294 597636 190350
rect 597704 190294 597760 190350
rect 597828 190294 597884 190350
rect 597456 190170 597512 190226
rect 597580 190170 597636 190226
rect 597704 190170 597760 190226
rect 597828 190170 597884 190226
rect 597456 190046 597512 190102
rect 597580 190046 597636 190102
rect 597704 190046 597760 190102
rect 597828 190046 597884 190102
rect 597456 189922 597512 189978
rect 597580 189922 597636 189978
rect 597704 189922 597760 189978
rect 597828 189922 597884 189978
rect 597456 172294 597512 172350
rect 597580 172294 597636 172350
rect 597704 172294 597760 172350
rect 597828 172294 597884 172350
rect 597456 172170 597512 172226
rect 597580 172170 597636 172226
rect 597704 172170 597760 172226
rect 597828 172170 597884 172226
rect 597456 172046 597512 172102
rect 597580 172046 597636 172102
rect 597704 172046 597760 172102
rect 597828 172046 597884 172102
rect 597456 171922 597512 171978
rect 597580 171922 597636 171978
rect 597704 171922 597760 171978
rect 597828 171922 597884 171978
rect 597456 154294 597512 154350
rect 597580 154294 597636 154350
rect 597704 154294 597760 154350
rect 597828 154294 597884 154350
rect 597456 154170 597512 154226
rect 597580 154170 597636 154226
rect 597704 154170 597760 154226
rect 597828 154170 597884 154226
rect 597456 154046 597512 154102
rect 597580 154046 597636 154102
rect 597704 154046 597760 154102
rect 597828 154046 597884 154102
rect 597456 153922 597512 153978
rect 597580 153922 597636 153978
rect 597704 153922 597760 153978
rect 597828 153922 597884 153978
rect 597456 136294 597512 136350
rect 597580 136294 597636 136350
rect 597704 136294 597760 136350
rect 597828 136294 597884 136350
rect 597456 136170 597512 136226
rect 597580 136170 597636 136226
rect 597704 136170 597760 136226
rect 597828 136170 597884 136226
rect 597456 136046 597512 136102
rect 597580 136046 597636 136102
rect 597704 136046 597760 136102
rect 597828 136046 597884 136102
rect 597456 135922 597512 135978
rect 597580 135922 597636 135978
rect 597704 135922 597760 135978
rect 597828 135922 597884 135978
rect 597456 118294 597512 118350
rect 597580 118294 597636 118350
rect 597704 118294 597760 118350
rect 597828 118294 597884 118350
rect 597456 118170 597512 118226
rect 597580 118170 597636 118226
rect 597704 118170 597760 118226
rect 597828 118170 597884 118226
rect 597456 118046 597512 118102
rect 597580 118046 597636 118102
rect 597704 118046 597760 118102
rect 597828 118046 597884 118102
rect 597456 117922 597512 117978
rect 597580 117922 597636 117978
rect 597704 117922 597760 117978
rect 597828 117922 597884 117978
rect 597456 100294 597512 100350
rect 597580 100294 597636 100350
rect 597704 100294 597760 100350
rect 597828 100294 597884 100350
rect 597456 100170 597512 100226
rect 597580 100170 597636 100226
rect 597704 100170 597760 100226
rect 597828 100170 597884 100226
rect 597456 100046 597512 100102
rect 597580 100046 597636 100102
rect 597704 100046 597760 100102
rect 597828 100046 597884 100102
rect 597456 99922 597512 99978
rect 597580 99922 597636 99978
rect 597704 99922 597760 99978
rect 597828 99922 597884 99978
rect 597456 82294 597512 82350
rect 597580 82294 597636 82350
rect 597704 82294 597760 82350
rect 597828 82294 597884 82350
rect 597456 82170 597512 82226
rect 597580 82170 597636 82226
rect 597704 82170 597760 82226
rect 597828 82170 597884 82226
rect 597456 82046 597512 82102
rect 597580 82046 597636 82102
rect 597704 82046 597760 82102
rect 597828 82046 597884 82102
rect 597456 81922 597512 81978
rect 597580 81922 597636 81978
rect 597704 81922 597760 81978
rect 597828 81922 597884 81978
rect 597456 64294 597512 64350
rect 597580 64294 597636 64350
rect 597704 64294 597760 64350
rect 597828 64294 597884 64350
rect 597456 64170 597512 64226
rect 597580 64170 597636 64226
rect 597704 64170 597760 64226
rect 597828 64170 597884 64226
rect 597456 64046 597512 64102
rect 597580 64046 597636 64102
rect 597704 64046 597760 64102
rect 597828 64046 597884 64102
rect 597456 63922 597512 63978
rect 597580 63922 597636 63978
rect 597704 63922 597760 63978
rect 597828 63922 597884 63978
rect 597456 46294 597512 46350
rect 597580 46294 597636 46350
rect 597704 46294 597760 46350
rect 597828 46294 597884 46350
rect 597456 46170 597512 46226
rect 597580 46170 597636 46226
rect 597704 46170 597760 46226
rect 597828 46170 597884 46226
rect 597456 46046 597512 46102
rect 597580 46046 597636 46102
rect 597704 46046 597760 46102
rect 597828 46046 597884 46102
rect 597456 45922 597512 45978
rect 597580 45922 597636 45978
rect 597704 45922 597760 45978
rect 597828 45922 597884 45978
rect 597456 28294 597512 28350
rect 597580 28294 597636 28350
rect 597704 28294 597760 28350
rect 597828 28294 597884 28350
rect 597456 28170 597512 28226
rect 597580 28170 597636 28226
rect 597704 28170 597760 28226
rect 597828 28170 597884 28226
rect 597456 28046 597512 28102
rect 597580 28046 597636 28102
rect 597704 28046 597760 28102
rect 597828 28046 597884 28102
rect 597456 27922 597512 27978
rect 597580 27922 597636 27978
rect 597704 27922 597760 27978
rect 597828 27922 597884 27978
rect 597456 10294 597512 10350
rect 597580 10294 597636 10350
rect 597704 10294 597760 10350
rect 597828 10294 597884 10350
rect 597456 10170 597512 10226
rect 597580 10170 597636 10226
rect 597704 10170 597760 10226
rect 597828 10170 597884 10226
rect 597456 10046 597512 10102
rect 597580 10046 597636 10102
rect 597704 10046 597760 10102
rect 597828 10046 597884 10102
rect 597456 9922 597512 9978
rect 597580 9922 597636 9978
rect 597704 9922 597760 9978
rect 597828 9922 597884 9978
rect 592914 -1176 592970 -1120
rect 593038 -1176 593094 -1120
rect 593162 -1176 593218 -1120
rect 593286 -1176 593342 -1120
rect 592914 -1300 592970 -1244
rect 593038 -1300 593094 -1244
rect 593162 -1300 593218 -1244
rect 593286 -1300 593342 -1244
rect 592914 -1424 592970 -1368
rect 593038 -1424 593094 -1368
rect 593162 -1424 593218 -1368
rect 593286 -1424 593342 -1368
rect 592914 -1548 592970 -1492
rect 593038 -1548 593094 -1492
rect 593162 -1548 593218 -1492
rect 593286 -1548 593342 -1492
rect 597456 -1176 597512 -1120
rect 597580 -1176 597636 -1120
rect 597704 -1176 597760 -1120
rect 597828 -1176 597884 -1120
rect 597456 -1300 597512 -1244
rect 597580 -1300 597636 -1244
rect 597704 -1300 597760 -1244
rect 597828 -1300 597884 -1244
rect 597456 -1424 597512 -1368
rect 597580 -1424 597636 -1368
rect 597704 -1424 597760 -1368
rect 597828 -1424 597884 -1368
rect 597456 -1548 597512 -1492
rect 597580 -1548 597636 -1492
rect 597704 -1548 597760 -1492
rect 597828 -1548 597884 -1492
<< metal5 >>
rect -1916 598172 597980 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 9234 598172
rect 9290 598116 9358 598172
rect 9414 598116 9482 598172
rect 9538 598116 9606 598172
rect 9662 598116 39954 598172
rect 40010 598116 40078 598172
rect 40134 598116 40202 598172
rect 40258 598116 40326 598172
rect 40382 598116 70674 598172
rect 70730 598116 70798 598172
rect 70854 598116 70922 598172
rect 70978 598116 71046 598172
rect 71102 598116 101394 598172
rect 101450 598116 101518 598172
rect 101574 598116 101642 598172
rect 101698 598116 101766 598172
rect 101822 598116 132114 598172
rect 132170 598116 132238 598172
rect 132294 598116 132362 598172
rect 132418 598116 132486 598172
rect 132542 598116 162834 598172
rect 162890 598116 162958 598172
rect 163014 598116 163082 598172
rect 163138 598116 163206 598172
rect 163262 598116 193554 598172
rect 193610 598116 193678 598172
rect 193734 598116 193802 598172
rect 193858 598116 193926 598172
rect 193982 598116 224274 598172
rect 224330 598116 224398 598172
rect 224454 598116 224522 598172
rect 224578 598116 224646 598172
rect 224702 598116 254994 598172
rect 255050 598116 255118 598172
rect 255174 598116 255242 598172
rect 255298 598116 255366 598172
rect 255422 598116 285714 598172
rect 285770 598116 285838 598172
rect 285894 598116 285962 598172
rect 286018 598116 286086 598172
rect 286142 598116 316434 598172
rect 316490 598116 316558 598172
rect 316614 598116 316682 598172
rect 316738 598116 316806 598172
rect 316862 598116 347154 598172
rect 347210 598116 347278 598172
rect 347334 598116 347402 598172
rect 347458 598116 347526 598172
rect 347582 598116 377874 598172
rect 377930 598116 377998 598172
rect 378054 598116 378122 598172
rect 378178 598116 378246 598172
rect 378302 598116 408594 598172
rect 408650 598116 408718 598172
rect 408774 598116 408842 598172
rect 408898 598116 408966 598172
rect 409022 598116 439314 598172
rect 439370 598116 439438 598172
rect 439494 598116 439562 598172
rect 439618 598116 439686 598172
rect 439742 598116 470034 598172
rect 470090 598116 470158 598172
rect 470214 598116 470282 598172
rect 470338 598116 470406 598172
rect 470462 598116 500754 598172
rect 500810 598116 500878 598172
rect 500934 598116 501002 598172
rect 501058 598116 501126 598172
rect 501182 598116 531474 598172
rect 531530 598116 531598 598172
rect 531654 598116 531722 598172
rect 531778 598116 531846 598172
rect 531902 598116 562194 598172
rect 562250 598116 562318 598172
rect 562374 598116 562442 598172
rect 562498 598116 562566 598172
rect 562622 598116 592914 598172
rect 592970 598116 593038 598172
rect 593094 598116 593162 598172
rect 593218 598116 593286 598172
rect 593342 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect -1916 598048 597980 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 9234 598048
rect 9290 597992 9358 598048
rect 9414 597992 9482 598048
rect 9538 597992 9606 598048
rect 9662 597992 39954 598048
rect 40010 597992 40078 598048
rect 40134 597992 40202 598048
rect 40258 597992 40326 598048
rect 40382 597992 70674 598048
rect 70730 597992 70798 598048
rect 70854 597992 70922 598048
rect 70978 597992 71046 598048
rect 71102 597992 101394 598048
rect 101450 597992 101518 598048
rect 101574 597992 101642 598048
rect 101698 597992 101766 598048
rect 101822 597992 132114 598048
rect 132170 597992 132238 598048
rect 132294 597992 132362 598048
rect 132418 597992 132486 598048
rect 132542 597992 162834 598048
rect 162890 597992 162958 598048
rect 163014 597992 163082 598048
rect 163138 597992 163206 598048
rect 163262 597992 193554 598048
rect 193610 597992 193678 598048
rect 193734 597992 193802 598048
rect 193858 597992 193926 598048
rect 193982 597992 224274 598048
rect 224330 597992 224398 598048
rect 224454 597992 224522 598048
rect 224578 597992 224646 598048
rect 224702 597992 254994 598048
rect 255050 597992 255118 598048
rect 255174 597992 255242 598048
rect 255298 597992 255366 598048
rect 255422 597992 285714 598048
rect 285770 597992 285838 598048
rect 285894 597992 285962 598048
rect 286018 597992 286086 598048
rect 286142 597992 316434 598048
rect 316490 597992 316558 598048
rect 316614 597992 316682 598048
rect 316738 597992 316806 598048
rect 316862 597992 347154 598048
rect 347210 597992 347278 598048
rect 347334 597992 347402 598048
rect 347458 597992 347526 598048
rect 347582 597992 377874 598048
rect 377930 597992 377998 598048
rect 378054 597992 378122 598048
rect 378178 597992 378246 598048
rect 378302 597992 408594 598048
rect 408650 597992 408718 598048
rect 408774 597992 408842 598048
rect 408898 597992 408966 598048
rect 409022 597992 439314 598048
rect 439370 597992 439438 598048
rect 439494 597992 439562 598048
rect 439618 597992 439686 598048
rect 439742 597992 470034 598048
rect 470090 597992 470158 598048
rect 470214 597992 470282 598048
rect 470338 597992 470406 598048
rect 470462 597992 500754 598048
rect 500810 597992 500878 598048
rect 500934 597992 501002 598048
rect 501058 597992 501126 598048
rect 501182 597992 531474 598048
rect 531530 597992 531598 598048
rect 531654 597992 531722 598048
rect 531778 597992 531846 598048
rect 531902 597992 562194 598048
rect 562250 597992 562318 598048
rect 562374 597992 562442 598048
rect 562498 597992 562566 598048
rect 562622 597992 592914 598048
rect 592970 597992 593038 598048
rect 593094 597992 593162 598048
rect 593218 597992 593286 598048
rect 593342 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect -1916 597924 597980 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 9234 597924
rect 9290 597868 9358 597924
rect 9414 597868 9482 597924
rect 9538 597868 9606 597924
rect 9662 597868 39954 597924
rect 40010 597868 40078 597924
rect 40134 597868 40202 597924
rect 40258 597868 40326 597924
rect 40382 597868 70674 597924
rect 70730 597868 70798 597924
rect 70854 597868 70922 597924
rect 70978 597868 71046 597924
rect 71102 597868 101394 597924
rect 101450 597868 101518 597924
rect 101574 597868 101642 597924
rect 101698 597868 101766 597924
rect 101822 597868 132114 597924
rect 132170 597868 132238 597924
rect 132294 597868 132362 597924
rect 132418 597868 132486 597924
rect 132542 597868 162834 597924
rect 162890 597868 162958 597924
rect 163014 597868 163082 597924
rect 163138 597868 163206 597924
rect 163262 597868 193554 597924
rect 193610 597868 193678 597924
rect 193734 597868 193802 597924
rect 193858 597868 193926 597924
rect 193982 597868 224274 597924
rect 224330 597868 224398 597924
rect 224454 597868 224522 597924
rect 224578 597868 224646 597924
rect 224702 597868 254994 597924
rect 255050 597868 255118 597924
rect 255174 597868 255242 597924
rect 255298 597868 255366 597924
rect 255422 597868 285714 597924
rect 285770 597868 285838 597924
rect 285894 597868 285962 597924
rect 286018 597868 286086 597924
rect 286142 597868 316434 597924
rect 316490 597868 316558 597924
rect 316614 597868 316682 597924
rect 316738 597868 316806 597924
rect 316862 597868 347154 597924
rect 347210 597868 347278 597924
rect 347334 597868 347402 597924
rect 347458 597868 347526 597924
rect 347582 597868 377874 597924
rect 377930 597868 377998 597924
rect 378054 597868 378122 597924
rect 378178 597868 378246 597924
rect 378302 597868 408594 597924
rect 408650 597868 408718 597924
rect 408774 597868 408842 597924
rect 408898 597868 408966 597924
rect 409022 597868 439314 597924
rect 439370 597868 439438 597924
rect 439494 597868 439562 597924
rect 439618 597868 439686 597924
rect 439742 597868 470034 597924
rect 470090 597868 470158 597924
rect 470214 597868 470282 597924
rect 470338 597868 470406 597924
rect 470462 597868 500754 597924
rect 500810 597868 500878 597924
rect 500934 597868 501002 597924
rect 501058 597868 501126 597924
rect 501182 597868 531474 597924
rect 531530 597868 531598 597924
rect 531654 597868 531722 597924
rect 531778 597868 531846 597924
rect 531902 597868 562194 597924
rect 562250 597868 562318 597924
rect 562374 597868 562442 597924
rect 562498 597868 562566 597924
rect 562622 597868 592914 597924
rect 592970 597868 593038 597924
rect 593094 597868 593162 597924
rect 593218 597868 593286 597924
rect 593342 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect -1916 597800 597980 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 9234 597800
rect 9290 597744 9358 597800
rect 9414 597744 9482 597800
rect 9538 597744 9606 597800
rect 9662 597744 39954 597800
rect 40010 597744 40078 597800
rect 40134 597744 40202 597800
rect 40258 597744 40326 597800
rect 40382 597744 70674 597800
rect 70730 597744 70798 597800
rect 70854 597744 70922 597800
rect 70978 597744 71046 597800
rect 71102 597744 101394 597800
rect 101450 597744 101518 597800
rect 101574 597744 101642 597800
rect 101698 597744 101766 597800
rect 101822 597744 132114 597800
rect 132170 597744 132238 597800
rect 132294 597744 132362 597800
rect 132418 597744 132486 597800
rect 132542 597744 162834 597800
rect 162890 597744 162958 597800
rect 163014 597744 163082 597800
rect 163138 597744 163206 597800
rect 163262 597744 193554 597800
rect 193610 597744 193678 597800
rect 193734 597744 193802 597800
rect 193858 597744 193926 597800
rect 193982 597744 224274 597800
rect 224330 597744 224398 597800
rect 224454 597744 224522 597800
rect 224578 597744 224646 597800
rect 224702 597744 254994 597800
rect 255050 597744 255118 597800
rect 255174 597744 255242 597800
rect 255298 597744 255366 597800
rect 255422 597744 285714 597800
rect 285770 597744 285838 597800
rect 285894 597744 285962 597800
rect 286018 597744 286086 597800
rect 286142 597744 316434 597800
rect 316490 597744 316558 597800
rect 316614 597744 316682 597800
rect 316738 597744 316806 597800
rect 316862 597744 347154 597800
rect 347210 597744 347278 597800
rect 347334 597744 347402 597800
rect 347458 597744 347526 597800
rect 347582 597744 377874 597800
rect 377930 597744 377998 597800
rect 378054 597744 378122 597800
rect 378178 597744 378246 597800
rect 378302 597744 408594 597800
rect 408650 597744 408718 597800
rect 408774 597744 408842 597800
rect 408898 597744 408966 597800
rect 409022 597744 439314 597800
rect 439370 597744 439438 597800
rect 439494 597744 439562 597800
rect 439618 597744 439686 597800
rect 439742 597744 470034 597800
rect 470090 597744 470158 597800
rect 470214 597744 470282 597800
rect 470338 597744 470406 597800
rect 470462 597744 500754 597800
rect 500810 597744 500878 597800
rect 500934 597744 501002 597800
rect 501058 597744 501126 597800
rect 501182 597744 531474 597800
rect 531530 597744 531598 597800
rect 531654 597744 531722 597800
rect 531778 597744 531846 597800
rect 531902 597744 562194 597800
rect 562250 597744 562318 597800
rect 562374 597744 562442 597800
rect 562498 597744 562566 597800
rect 562622 597744 592914 597800
rect 592970 597744 593038 597800
rect 593094 597744 593162 597800
rect 593218 597744 593286 597800
rect 593342 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect -1916 597648 597980 597744
rect -956 597212 597020 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 5514 597212
rect 5570 597156 5638 597212
rect 5694 597156 5762 597212
rect 5818 597156 5886 597212
rect 5942 597156 589194 597212
rect 589250 597156 589318 597212
rect 589374 597156 589442 597212
rect 589498 597156 589566 597212
rect 589622 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect -956 597088 597020 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 5514 597088
rect 5570 597032 5638 597088
rect 5694 597032 5762 597088
rect 5818 597032 5886 597088
rect 5942 597032 589194 597088
rect 589250 597032 589318 597088
rect 589374 597032 589442 597088
rect 589498 597032 589566 597088
rect 589622 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect -956 596964 597020 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 5514 596964
rect 5570 596908 5638 596964
rect 5694 596908 5762 596964
rect 5818 596908 5886 596964
rect 5942 596908 589194 596964
rect 589250 596908 589318 596964
rect 589374 596908 589442 596964
rect 589498 596908 589566 596964
rect 589622 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect -956 596840 597020 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 5514 596840
rect 5570 596784 5638 596840
rect 5694 596784 5762 596840
rect 5818 596784 5886 596840
rect 5942 596784 589194 596840
rect 589250 596784 589318 596840
rect 589374 596784 589442 596840
rect 589498 596784 589566 596840
rect 589622 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect -956 596688 597020 596784
rect -1916 586350 597980 586446
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 9234 586350
rect 9290 586294 9358 586350
rect 9414 586294 9482 586350
rect 9538 586294 9606 586350
rect 9662 586294 39954 586350
rect 40010 586294 40078 586350
rect 40134 586294 40202 586350
rect 40258 586294 40326 586350
rect 40382 586294 70674 586350
rect 70730 586294 70798 586350
rect 70854 586294 70922 586350
rect 70978 586294 71046 586350
rect 71102 586294 101394 586350
rect 101450 586294 101518 586350
rect 101574 586294 101642 586350
rect 101698 586294 101766 586350
rect 101822 586294 132114 586350
rect 132170 586294 132238 586350
rect 132294 586294 132362 586350
rect 132418 586294 132486 586350
rect 132542 586294 162834 586350
rect 162890 586294 162958 586350
rect 163014 586294 163082 586350
rect 163138 586294 163206 586350
rect 163262 586294 193554 586350
rect 193610 586294 193678 586350
rect 193734 586294 193802 586350
rect 193858 586294 193926 586350
rect 193982 586294 224274 586350
rect 224330 586294 224398 586350
rect 224454 586294 224522 586350
rect 224578 586294 224646 586350
rect 224702 586294 254994 586350
rect 255050 586294 255118 586350
rect 255174 586294 255242 586350
rect 255298 586294 255366 586350
rect 255422 586294 285714 586350
rect 285770 586294 285838 586350
rect 285894 586294 285962 586350
rect 286018 586294 286086 586350
rect 286142 586294 316434 586350
rect 316490 586294 316558 586350
rect 316614 586294 316682 586350
rect 316738 586294 316806 586350
rect 316862 586294 347154 586350
rect 347210 586294 347278 586350
rect 347334 586294 347402 586350
rect 347458 586294 347526 586350
rect 347582 586294 377874 586350
rect 377930 586294 377998 586350
rect 378054 586294 378122 586350
rect 378178 586294 378246 586350
rect 378302 586294 408594 586350
rect 408650 586294 408718 586350
rect 408774 586294 408842 586350
rect 408898 586294 408966 586350
rect 409022 586294 439314 586350
rect 439370 586294 439438 586350
rect 439494 586294 439562 586350
rect 439618 586294 439686 586350
rect 439742 586294 470034 586350
rect 470090 586294 470158 586350
rect 470214 586294 470282 586350
rect 470338 586294 470406 586350
rect 470462 586294 500754 586350
rect 500810 586294 500878 586350
rect 500934 586294 501002 586350
rect 501058 586294 501126 586350
rect 501182 586294 531474 586350
rect 531530 586294 531598 586350
rect 531654 586294 531722 586350
rect 531778 586294 531846 586350
rect 531902 586294 562194 586350
rect 562250 586294 562318 586350
rect 562374 586294 562442 586350
rect 562498 586294 562566 586350
rect 562622 586294 592914 586350
rect 592970 586294 593038 586350
rect 593094 586294 593162 586350
rect 593218 586294 593286 586350
rect 593342 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect -1916 586226 597980 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 9234 586226
rect 9290 586170 9358 586226
rect 9414 586170 9482 586226
rect 9538 586170 9606 586226
rect 9662 586170 39954 586226
rect 40010 586170 40078 586226
rect 40134 586170 40202 586226
rect 40258 586170 40326 586226
rect 40382 586170 70674 586226
rect 70730 586170 70798 586226
rect 70854 586170 70922 586226
rect 70978 586170 71046 586226
rect 71102 586170 101394 586226
rect 101450 586170 101518 586226
rect 101574 586170 101642 586226
rect 101698 586170 101766 586226
rect 101822 586170 132114 586226
rect 132170 586170 132238 586226
rect 132294 586170 132362 586226
rect 132418 586170 132486 586226
rect 132542 586170 162834 586226
rect 162890 586170 162958 586226
rect 163014 586170 163082 586226
rect 163138 586170 163206 586226
rect 163262 586170 193554 586226
rect 193610 586170 193678 586226
rect 193734 586170 193802 586226
rect 193858 586170 193926 586226
rect 193982 586170 224274 586226
rect 224330 586170 224398 586226
rect 224454 586170 224522 586226
rect 224578 586170 224646 586226
rect 224702 586170 254994 586226
rect 255050 586170 255118 586226
rect 255174 586170 255242 586226
rect 255298 586170 255366 586226
rect 255422 586170 285714 586226
rect 285770 586170 285838 586226
rect 285894 586170 285962 586226
rect 286018 586170 286086 586226
rect 286142 586170 316434 586226
rect 316490 586170 316558 586226
rect 316614 586170 316682 586226
rect 316738 586170 316806 586226
rect 316862 586170 347154 586226
rect 347210 586170 347278 586226
rect 347334 586170 347402 586226
rect 347458 586170 347526 586226
rect 347582 586170 377874 586226
rect 377930 586170 377998 586226
rect 378054 586170 378122 586226
rect 378178 586170 378246 586226
rect 378302 586170 408594 586226
rect 408650 586170 408718 586226
rect 408774 586170 408842 586226
rect 408898 586170 408966 586226
rect 409022 586170 439314 586226
rect 439370 586170 439438 586226
rect 439494 586170 439562 586226
rect 439618 586170 439686 586226
rect 439742 586170 470034 586226
rect 470090 586170 470158 586226
rect 470214 586170 470282 586226
rect 470338 586170 470406 586226
rect 470462 586170 500754 586226
rect 500810 586170 500878 586226
rect 500934 586170 501002 586226
rect 501058 586170 501126 586226
rect 501182 586170 531474 586226
rect 531530 586170 531598 586226
rect 531654 586170 531722 586226
rect 531778 586170 531846 586226
rect 531902 586170 562194 586226
rect 562250 586170 562318 586226
rect 562374 586170 562442 586226
rect 562498 586170 562566 586226
rect 562622 586170 592914 586226
rect 592970 586170 593038 586226
rect 593094 586170 593162 586226
rect 593218 586170 593286 586226
rect 593342 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect -1916 586102 597980 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 9234 586102
rect 9290 586046 9358 586102
rect 9414 586046 9482 586102
rect 9538 586046 9606 586102
rect 9662 586046 39954 586102
rect 40010 586046 40078 586102
rect 40134 586046 40202 586102
rect 40258 586046 40326 586102
rect 40382 586046 70674 586102
rect 70730 586046 70798 586102
rect 70854 586046 70922 586102
rect 70978 586046 71046 586102
rect 71102 586046 101394 586102
rect 101450 586046 101518 586102
rect 101574 586046 101642 586102
rect 101698 586046 101766 586102
rect 101822 586046 132114 586102
rect 132170 586046 132238 586102
rect 132294 586046 132362 586102
rect 132418 586046 132486 586102
rect 132542 586046 162834 586102
rect 162890 586046 162958 586102
rect 163014 586046 163082 586102
rect 163138 586046 163206 586102
rect 163262 586046 193554 586102
rect 193610 586046 193678 586102
rect 193734 586046 193802 586102
rect 193858 586046 193926 586102
rect 193982 586046 224274 586102
rect 224330 586046 224398 586102
rect 224454 586046 224522 586102
rect 224578 586046 224646 586102
rect 224702 586046 254994 586102
rect 255050 586046 255118 586102
rect 255174 586046 255242 586102
rect 255298 586046 255366 586102
rect 255422 586046 285714 586102
rect 285770 586046 285838 586102
rect 285894 586046 285962 586102
rect 286018 586046 286086 586102
rect 286142 586046 316434 586102
rect 316490 586046 316558 586102
rect 316614 586046 316682 586102
rect 316738 586046 316806 586102
rect 316862 586046 347154 586102
rect 347210 586046 347278 586102
rect 347334 586046 347402 586102
rect 347458 586046 347526 586102
rect 347582 586046 377874 586102
rect 377930 586046 377998 586102
rect 378054 586046 378122 586102
rect 378178 586046 378246 586102
rect 378302 586046 408594 586102
rect 408650 586046 408718 586102
rect 408774 586046 408842 586102
rect 408898 586046 408966 586102
rect 409022 586046 439314 586102
rect 439370 586046 439438 586102
rect 439494 586046 439562 586102
rect 439618 586046 439686 586102
rect 439742 586046 470034 586102
rect 470090 586046 470158 586102
rect 470214 586046 470282 586102
rect 470338 586046 470406 586102
rect 470462 586046 500754 586102
rect 500810 586046 500878 586102
rect 500934 586046 501002 586102
rect 501058 586046 501126 586102
rect 501182 586046 531474 586102
rect 531530 586046 531598 586102
rect 531654 586046 531722 586102
rect 531778 586046 531846 586102
rect 531902 586046 562194 586102
rect 562250 586046 562318 586102
rect 562374 586046 562442 586102
rect 562498 586046 562566 586102
rect 562622 586046 592914 586102
rect 592970 586046 593038 586102
rect 593094 586046 593162 586102
rect 593218 586046 593286 586102
rect 593342 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect -1916 585978 597980 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 9234 585978
rect 9290 585922 9358 585978
rect 9414 585922 9482 585978
rect 9538 585922 9606 585978
rect 9662 585922 39954 585978
rect 40010 585922 40078 585978
rect 40134 585922 40202 585978
rect 40258 585922 40326 585978
rect 40382 585922 70674 585978
rect 70730 585922 70798 585978
rect 70854 585922 70922 585978
rect 70978 585922 71046 585978
rect 71102 585922 101394 585978
rect 101450 585922 101518 585978
rect 101574 585922 101642 585978
rect 101698 585922 101766 585978
rect 101822 585922 132114 585978
rect 132170 585922 132238 585978
rect 132294 585922 132362 585978
rect 132418 585922 132486 585978
rect 132542 585922 162834 585978
rect 162890 585922 162958 585978
rect 163014 585922 163082 585978
rect 163138 585922 163206 585978
rect 163262 585922 193554 585978
rect 193610 585922 193678 585978
rect 193734 585922 193802 585978
rect 193858 585922 193926 585978
rect 193982 585922 224274 585978
rect 224330 585922 224398 585978
rect 224454 585922 224522 585978
rect 224578 585922 224646 585978
rect 224702 585922 254994 585978
rect 255050 585922 255118 585978
rect 255174 585922 255242 585978
rect 255298 585922 255366 585978
rect 255422 585922 285714 585978
rect 285770 585922 285838 585978
rect 285894 585922 285962 585978
rect 286018 585922 286086 585978
rect 286142 585922 316434 585978
rect 316490 585922 316558 585978
rect 316614 585922 316682 585978
rect 316738 585922 316806 585978
rect 316862 585922 347154 585978
rect 347210 585922 347278 585978
rect 347334 585922 347402 585978
rect 347458 585922 347526 585978
rect 347582 585922 377874 585978
rect 377930 585922 377998 585978
rect 378054 585922 378122 585978
rect 378178 585922 378246 585978
rect 378302 585922 408594 585978
rect 408650 585922 408718 585978
rect 408774 585922 408842 585978
rect 408898 585922 408966 585978
rect 409022 585922 439314 585978
rect 439370 585922 439438 585978
rect 439494 585922 439562 585978
rect 439618 585922 439686 585978
rect 439742 585922 470034 585978
rect 470090 585922 470158 585978
rect 470214 585922 470282 585978
rect 470338 585922 470406 585978
rect 470462 585922 500754 585978
rect 500810 585922 500878 585978
rect 500934 585922 501002 585978
rect 501058 585922 501126 585978
rect 501182 585922 531474 585978
rect 531530 585922 531598 585978
rect 531654 585922 531722 585978
rect 531778 585922 531846 585978
rect 531902 585922 562194 585978
rect 562250 585922 562318 585978
rect 562374 585922 562442 585978
rect 562498 585922 562566 585978
rect 562622 585922 592914 585978
rect 592970 585922 593038 585978
rect 593094 585922 593162 585978
rect 593218 585922 593286 585978
rect 593342 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect -1916 585826 597980 585922
rect -1916 580350 597980 580446
rect -1916 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 5514 580350
rect 5570 580294 5638 580350
rect 5694 580294 5762 580350
rect 5818 580294 5886 580350
rect 5942 580294 12518 580350
rect 12574 580294 12642 580350
rect 12698 580294 43238 580350
rect 43294 580294 43362 580350
rect 43418 580294 73958 580350
rect 74014 580294 74082 580350
rect 74138 580294 104678 580350
rect 104734 580294 104802 580350
rect 104858 580294 135398 580350
rect 135454 580294 135522 580350
rect 135578 580294 166118 580350
rect 166174 580294 166242 580350
rect 166298 580294 196838 580350
rect 196894 580294 196962 580350
rect 197018 580294 227558 580350
rect 227614 580294 227682 580350
rect 227738 580294 258278 580350
rect 258334 580294 258402 580350
rect 258458 580294 288998 580350
rect 289054 580294 289122 580350
rect 289178 580294 319718 580350
rect 319774 580294 319842 580350
rect 319898 580294 350438 580350
rect 350494 580294 350562 580350
rect 350618 580294 381158 580350
rect 381214 580294 381282 580350
rect 381338 580294 411878 580350
rect 411934 580294 412002 580350
rect 412058 580294 442598 580350
rect 442654 580294 442722 580350
rect 442778 580294 473318 580350
rect 473374 580294 473442 580350
rect 473498 580294 504038 580350
rect 504094 580294 504162 580350
rect 504218 580294 534758 580350
rect 534814 580294 534882 580350
rect 534938 580294 565478 580350
rect 565534 580294 565602 580350
rect 565658 580294 589194 580350
rect 589250 580294 589318 580350
rect 589374 580294 589442 580350
rect 589498 580294 589566 580350
rect 589622 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597980 580350
rect -1916 580226 597980 580294
rect -1916 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 5514 580226
rect 5570 580170 5638 580226
rect 5694 580170 5762 580226
rect 5818 580170 5886 580226
rect 5942 580170 12518 580226
rect 12574 580170 12642 580226
rect 12698 580170 43238 580226
rect 43294 580170 43362 580226
rect 43418 580170 73958 580226
rect 74014 580170 74082 580226
rect 74138 580170 104678 580226
rect 104734 580170 104802 580226
rect 104858 580170 135398 580226
rect 135454 580170 135522 580226
rect 135578 580170 166118 580226
rect 166174 580170 166242 580226
rect 166298 580170 196838 580226
rect 196894 580170 196962 580226
rect 197018 580170 227558 580226
rect 227614 580170 227682 580226
rect 227738 580170 258278 580226
rect 258334 580170 258402 580226
rect 258458 580170 288998 580226
rect 289054 580170 289122 580226
rect 289178 580170 319718 580226
rect 319774 580170 319842 580226
rect 319898 580170 350438 580226
rect 350494 580170 350562 580226
rect 350618 580170 381158 580226
rect 381214 580170 381282 580226
rect 381338 580170 411878 580226
rect 411934 580170 412002 580226
rect 412058 580170 442598 580226
rect 442654 580170 442722 580226
rect 442778 580170 473318 580226
rect 473374 580170 473442 580226
rect 473498 580170 504038 580226
rect 504094 580170 504162 580226
rect 504218 580170 534758 580226
rect 534814 580170 534882 580226
rect 534938 580170 565478 580226
rect 565534 580170 565602 580226
rect 565658 580170 589194 580226
rect 589250 580170 589318 580226
rect 589374 580170 589442 580226
rect 589498 580170 589566 580226
rect 589622 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597980 580226
rect -1916 580102 597980 580170
rect -1916 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 5514 580102
rect 5570 580046 5638 580102
rect 5694 580046 5762 580102
rect 5818 580046 5886 580102
rect 5942 580046 12518 580102
rect 12574 580046 12642 580102
rect 12698 580046 43238 580102
rect 43294 580046 43362 580102
rect 43418 580046 73958 580102
rect 74014 580046 74082 580102
rect 74138 580046 104678 580102
rect 104734 580046 104802 580102
rect 104858 580046 135398 580102
rect 135454 580046 135522 580102
rect 135578 580046 166118 580102
rect 166174 580046 166242 580102
rect 166298 580046 196838 580102
rect 196894 580046 196962 580102
rect 197018 580046 227558 580102
rect 227614 580046 227682 580102
rect 227738 580046 258278 580102
rect 258334 580046 258402 580102
rect 258458 580046 288998 580102
rect 289054 580046 289122 580102
rect 289178 580046 319718 580102
rect 319774 580046 319842 580102
rect 319898 580046 350438 580102
rect 350494 580046 350562 580102
rect 350618 580046 381158 580102
rect 381214 580046 381282 580102
rect 381338 580046 411878 580102
rect 411934 580046 412002 580102
rect 412058 580046 442598 580102
rect 442654 580046 442722 580102
rect 442778 580046 473318 580102
rect 473374 580046 473442 580102
rect 473498 580046 504038 580102
rect 504094 580046 504162 580102
rect 504218 580046 534758 580102
rect 534814 580046 534882 580102
rect 534938 580046 565478 580102
rect 565534 580046 565602 580102
rect 565658 580046 589194 580102
rect 589250 580046 589318 580102
rect 589374 580046 589442 580102
rect 589498 580046 589566 580102
rect 589622 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597980 580102
rect -1916 579978 597980 580046
rect -1916 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 5514 579978
rect 5570 579922 5638 579978
rect 5694 579922 5762 579978
rect 5818 579922 5886 579978
rect 5942 579922 12518 579978
rect 12574 579922 12642 579978
rect 12698 579922 43238 579978
rect 43294 579922 43362 579978
rect 43418 579922 73958 579978
rect 74014 579922 74082 579978
rect 74138 579922 104678 579978
rect 104734 579922 104802 579978
rect 104858 579922 135398 579978
rect 135454 579922 135522 579978
rect 135578 579922 166118 579978
rect 166174 579922 166242 579978
rect 166298 579922 196838 579978
rect 196894 579922 196962 579978
rect 197018 579922 227558 579978
rect 227614 579922 227682 579978
rect 227738 579922 258278 579978
rect 258334 579922 258402 579978
rect 258458 579922 288998 579978
rect 289054 579922 289122 579978
rect 289178 579922 319718 579978
rect 319774 579922 319842 579978
rect 319898 579922 350438 579978
rect 350494 579922 350562 579978
rect 350618 579922 381158 579978
rect 381214 579922 381282 579978
rect 381338 579922 411878 579978
rect 411934 579922 412002 579978
rect 412058 579922 442598 579978
rect 442654 579922 442722 579978
rect 442778 579922 473318 579978
rect 473374 579922 473442 579978
rect 473498 579922 504038 579978
rect 504094 579922 504162 579978
rect 504218 579922 534758 579978
rect 534814 579922 534882 579978
rect 534938 579922 565478 579978
rect 565534 579922 565602 579978
rect 565658 579922 589194 579978
rect 589250 579922 589318 579978
rect 589374 579922 589442 579978
rect 589498 579922 589566 579978
rect 589622 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597980 579978
rect -1916 579826 597980 579922
rect -1916 568350 597980 568446
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 27878 568350
rect 27934 568294 28002 568350
rect 28058 568294 58598 568350
rect 58654 568294 58722 568350
rect 58778 568294 89318 568350
rect 89374 568294 89442 568350
rect 89498 568294 120038 568350
rect 120094 568294 120162 568350
rect 120218 568294 150758 568350
rect 150814 568294 150882 568350
rect 150938 568294 181478 568350
rect 181534 568294 181602 568350
rect 181658 568294 212198 568350
rect 212254 568294 212322 568350
rect 212378 568294 242918 568350
rect 242974 568294 243042 568350
rect 243098 568294 273638 568350
rect 273694 568294 273762 568350
rect 273818 568294 304358 568350
rect 304414 568294 304482 568350
rect 304538 568294 335078 568350
rect 335134 568294 335202 568350
rect 335258 568294 365798 568350
rect 365854 568294 365922 568350
rect 365978 568294 396518 568350
rect 396574 568294 396642 568350
rect 396698 568294 427238 568350
rect 427294 568294 427362 568350
rect 427418 568294 457958 568350
rect 458014 568294 458082 568350
rect 458138 568294 488678 568350
rect 488734 568294 488802 568350
rect 488858 568294 519398 568350
rect 519454 568294 519522 568350
rect 519578 568294 550118 568350
rect 550174 568294 550242 568350
rect 550298 568294 592914 568350
rect 592970 568294 593038 568350
rect 593094 568294 593162 568350
rect 593218 568294 593286 568350
rect 593342 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect -1916 568226 597980 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 27878 568226
rect 27934 568170 28002 568226
rect 28058 568170 58598 568226
rect 58654 568170 58722 568226
rect 58778 568170 89318 568226
rect 89374 568170 89442 568226
rect 89498 568170 120038 568226
rect 120094 568170 120162 568226
rect 120218 568170 150758 568226
rect 150814 568170 150882 568226
rect 150938 568170 181478 568226
rect 181534 568170 181602 568226
rect 181658 568170 212198 568226
rect 212254 568170 212322 568226
rect 212378 568170 242918 568226
rect 242974 568170 243042 568226
rect 243098 568170 273638 568226
rect 273694 568170 273762 568226
rect 273818 568170 304358 568226
rect 304414 568170 304482 568226
rect 304538 568170 335078 568226
rect 335134 568170 335202 568226
rect 335258 568170 365798 568226
rect 365854 568170 365922 568226
rect 365978 568170 396518 568226
rect 396574 568170 396642 568226
rect 396698 568170 427238 568226
rect 427294 568170 427362 568226
rect 427418 568170 457958 568226
rect 458014 568170 458082 568226
rect 458138 568170 488678 568226
rect 488734 568170 488802 568226
rect 488858 568170 519398 568226
rect 519454 568170 519522 568226
rect 519578 568170 550118 568226
rect 550174 568170 550242 568226
rect 550298 568170 592914 568226
rect 592970 568170 593038 568226
rect 593094 568170 593162 568226
rect 593218 568170 593286 568226
rect 593342 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect -1916 568102 597980 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 27878 568102
rect 27934 568046 28002 568102
rect 28058 568046 58598 568102
rect 58654 568046 58722 568102
rect 58778 568046 89318 568102
rect 89374 568046 89442 568102
rect 89498 568046 120038 568102
rect 120094 568046 120162 568102
rect 120218 568046 150758 568102
rect 150814 568046 150882 568102
rect 150938 568046 181478 568102
rect 181534 568046 181602 568102
rect 181658 568046 212198 568102
rect 212254 568046 212322 568102
rect 212378 568046 242918 568102
rect 242974 568046 243042 568102
rect 243098 568046 273638 568102
rect 273694 568046 273762 568102
rect 273818 568046 304358 568102
rect 304414 568046 304482 568102
rect 304538 568046 335078 568102
rect 335134 568046 335202 568102
rect 335258 568046 365798 568102
rect 365854 568046 365922 568102
rect 365978 568046 396518 568102
rect 396574 568046 396642 568102
rect 396698 568046 427238 568102
rect 427294 568046 427362 568102
rect 427418 568046 457958 568102
rect 458014 568046 458082 568102
rect 458138 568046 488678 568102
rect 488734 568046 488802 568102
rect 488858 568046 519398 568102
rect 519454 568046 519522 568102
rect 519578 568046 550118 568102
rect 550174 568046 550242 568102
rect 550298 568046 592914 568102
rect 592970 568046 593038 568102
rect 593094 568046 593162 568102
rect 593218 568046 593286 568102
rect 593342 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect -1916 567978 597980 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 27878 567978
rect 27934 567922 28002 567978
rect 28058 567922 58598 567978
rect 58654 567922 58722 567978
rect 58778 567922 89318 567978
rect 89374 567922 89442 567978
rect 89498 567922 120038 567978
rect 120094 567922 120162 567978
rect 120218 567922 150758 567978
rect 150814 567922 150882 567978
rect 150938 567922 181478 567978
rect 181534 567922 181602 567978
rect 181658 567922 212198 567978
rect 212254 567922 212322 567978
rect 212378 567922 242918 567978
rect 242974 567922 243042 567978
rect 243098 567922 273638 567978
rect 273694 567922 273762 567978
rect 273818 567922 304358 567978
rect 304414 567922 304482 567978
rect 304538 567922 335078 567978
rect 335134 567922 335202 567978
rect 335258 567922 365798 567978
rect 365854 567922 365922 567978
rect 365978 567922 396518 567978
rect 396574 567922 396642 567978
rect 396698 567922 427238 567978
rect 427294 567922 427362 567978
rect 427418 567922 457958 567978
rect 458014 567922 458082 567978
rect 458138 567922 488678 567978
rect 488734 567922 488802 567978
rect 488858 567922 519398 567978
rect 519454 567922 519522 567978
rect 519578 567922 550118 567978
rect 550174 567922 550242 567978
rect 550298 567922 592914 567978
rect 592970 567922 593038 567978
rect 593094 567922 593162 567978
rect 593218 567922 593286 567978
rect 593342 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect -1916 567826 597980 567922
rect -1916 562350 597980 562446
rect -1916 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 5514 562350
rect 5570 562294 5638 562350
rect 5694 562294 5762 562350
rect 5818 562294 5886 562350
rect 5942 562294 12518 562350
rect 12574 562294 12642 562350
rect 12698 562294 43238 562350
rect 43294 562294 43362 562350
rect 43418 562294 73958 562350
rect 74014 562294 74082 562350
rect 74138 562294 104678 562350
rect 104734 562294 104802 562350
rect 104858 562294 135398 562350
rect 135454 562294 135522 562350
rect 135578 562294 166118 562350
rect 166174 562294 166242 562350
rect 166298 562294 196838 562350
rect 196894 562294 196962 562350
rect 197018 562294 227558 562350
rect 227614 562294 227682 562350
rect 227738 562294 258278 562350
rect 258334 562294 258402 562350
rect 258458 562294 288998 562350
rect 289054 562294 289122 562350
rect 289178 562294 319718 562350
rect 319774 562294 319842 562350
rect 319898 562294 350438 562350
rect 350494 562294 350562 562350
rect 350618 562294 381158 562350
rect 381214 562294 381282 562350
rect 381338 562294 411878 562350
rect 411934 562294 412002 562350
rect 412058 562294 442598 562350
rect 442654 562294 442722 562350
rect 442778 562294 473318 562350
rect 473374 562294 473442 562350
rect 473498 562294 504038 562350
rect 504094 562294 504162 562350
rect 504218 562294 534758 562350
rect 534814 562294 534882 562350
rect 534938 562294 565478 562350
rect 565534 562294 565602 562350
rect 565658 562294 589194 562350
rect 589250 562294 589318 562350
rect 589374 562294 589442 562350
rect 589498 562294 589566 562350
rect 589622 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597980 562350
rect -1916 562226 597980 562294
rect -1916 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 5514 562226
rect 5570 562170 5638 562226
rect 5694 562170 5762 562226
rect 5818 562170 5886 562226
rect 5942 562170 12518 562226
rect 12574 562170 12642 562226
rect 12698 562170 43238 562226
rect 43294 562170 43362 562226
rect 43418 562170 73958 562226
rect 74014 562170 74082 562226
rect 74138 562170 104678 562226
rect 104734 562170 104802 562226
rect 104858 562170 135398 562226
rect 135454 562170 135522 562226
rect 135578 562170 166118 562226
rect 166174 562170 166242 562226
rect 166298 562170 196838 562226
rect 196894 562170 196962 562226
rect 197018 562170 227558 562226
rect 227614 562170 227682 562226
rect 227738 562170 258278 562226
rect 258334 562170 258402 562226
rect 258458 562170 288998 562226
rect 289054 562170 289122 562226
rect 289178 562170 319718 562226
rect 319774 562170 319842 562226
rect 319898 562170 350438 562226
rect 350494 562170 350562 562226
rect 350618 562170 381158 562226
rect 381214 562170 381282 562226
rect 381338 562170 411878 562226
rect 411934 562170 412002 562226
rect 412058 562170 442598 562226
rect 442654 562170 442722 562226
rect 442778 562170 473318 562226
rect 473374 562170 473442 562226
rect 473498 562170 504038 562226
rect 504094 562170 504162 562226
rect 504218 562170 534758 562226
rect 534814 562170 534882 562226
rect 534938 562170 565478 562226
rect 565534 562170 565602 562226
rect 565658 562170 589194 562226
rect 589250 562170 589318 562226
rect 589374 562170 589442 562226
rect 589498 562170 589566 562226
rect 589622 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597980 562226
rect -1916 562102 597980 562170
rect -1916 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 5514 562102
rect 5570 562046 5638 562102
rect 5694 562046 5762 562102
rect 5818 562046 5886 562102
rect 5942 562046 12518 562102
rect 12574 562046 12642 562102
rect 12698 562046 43238 562102
rect 43294 562046 43362 562102
rect 43418 562046 73958 562102
rect 74014 562046 74082 562102
rect 74138 562046 104678 562102
rect 104734 562046 104802 562102
rect 104858 562046 135398 562102
rect 135454 562046 135522 562102
rect 135578 562046 166118 562102
rect 166174 562046 166242 562102
rect 166298 562046 196838 562102
rect 196894 562046 196962 562102
rect 197018 562046 227558 562102
rect 227614 562046 227682 562102
rect 227738 562046 258278 562102
rect 258334 562046 258402 562102
rect 258458 562046 288998 562102
rect 289054 562046 289122 562102
rect 289178 562046 319718 562102
rect 319774 562046 319842 562102
rect 319898 562046 350438 562102
rect 350494 562046 350562 562102
rect 350618 562046 381158 562102
rect 381214 562046 381282 562102
rect 381338 562046 411878 562102
rect 411934 562046 412002 562102
rect 412058 562046 442598 562102
rect 442654 562046 442722 562102
rect 442778 562046 473318 562102
rect 473374 562046 473442 562102
rect 473498 562046 504038 562102
rect 504094 562046 504162 562102
rect 504218 562046 534758 562102
rect 534814 562046 534882 562102
rect 534938 562046 565478 562102
rect 565534 562046 565602 562102
rect 565658 562046 589194 562102
rect 589250 562046 589318 562102
rect 589374 562046 589442 562102
rect 589498 562046 589566 562102
rect 589622 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597980 562102
rect -1916 561978 597980 562046
rect -1916 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 5514 561978
rect 5570 561922 5638 561978
rect 5694 561922 5762 561978
rect 5818 561922 5886 561978
rect 5942 561922 12518 561978
rect 12574 561922 12642 561978
rect 12698 561922 43238 561978
rect 43294 561922 43362 561978
rect 43418 561922 73958 561978
rect 74014 561922 74082 561978
rect 74138 561922 104678 561978
rect 104734 561922 104802 561978
rect 104858 561922 135398 561978
rect 135454 561922 135522 561978
rect 135578 561922 166118 561978
rect 166174 561922 166242 561978
rect 166298 561922 196838 561978
rect 196894 561922 196962 561978
rect 197018 561922 227558 561978
rect 227614 561922 227682 561978
rect 227738 561922 258278 561978
rect 258334 561922 258402 561978
rect 258458 561922 288998 561978
rect 289054 561922 289122 561978
rect 289178 561922 319718 561978
rect 319774 561922 319842 561978
rect 319898 561922 350438 561978
rect 350494 561922 350562 561978
rect 350618 561922 381158 561978
rect 381214 561922 381282 561978
rect 381338 561922 411878 561978
rect 411934 561922 412002 561978
rect 412058 561922 442598 561978
rect 442654 561922 442722 561978
rect 442778 561922 473318 561978
rect 473374 561922 473442 561978
rect 473498 561922 504038 561978
rect 504094 561922 504162 561978
rect 504218 561922 534758 561978
rect 534814 561922 534882 561978
rect 534938 561922 565478 561978
rect 565534 561922 565602 561978
rect 565658 561922 589194 561978
rect 589250 561922 589318 561978
rect 589374 561922 589442 561978
rect 589498 561922 589566 561978
rect 589622 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597980 561978
rect -1916 561826 597980 561922
rect -1916 550350 597980 550446
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 27878 550350
rect 27934 550294 28002 550350
rect 28058 550294 58598 550350
rect 58654 550294 58722 550350
rect 58778 550294 89318 550350
rect 89374 550294 89442 550350
rect 89498 550294 120038 550350
rect 120094 550294 120162 550350
rect 120218 550294 150758 550350
rect 150814 550294 150882 550350
rect 150938 550294 181478 550350
rect 181534 550294 181602 550350
rect 181658 550294 212198 550350
rect 212254 550294 212322 550350
rect 212378 550294 242918 550350
rect 242974 550294 243042 550350
rect 243098 550294 273638 550350
rect 273694 550294 273762 550350
rect 273818 550294 304358 550350
rect 304414 550294 304482 550350
rect 304538 550294 335078 550350
rect 335134 550294 335202 550350
rect 335258 550294 365798 550350
rect 365854 550294 365922 550350
rect 365978 550294 396518 550350
rect 396574 550294 396642 550350
rect 396698 550294 427238 550350
rect 427294 550294 427362 550350
rect 427418 550294 457958 550350
rect 458014 550294 458082 550350
rect 458138 550294 488678 550350
rect 488734 550294 488802 550350
rect 488858 550294 519398 550350
rect 519454 550294 519522 550350
rect 519578 550294 550118 550350
rect 550174 550294 550242 550350
rect 550298 550294 592914 550350
rect 592970 550294 593038 550350
rect 593094 550294 593162 550350
rect 593218 550294 593286 550350
rect 593342 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect -1916 550226 597980 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 27878 550226
rect 27934 550170 28002 550226
rect 28058 550170 58598 550226
rect 58654 550170 58722 550226
rect 58778 550170 89318 550226
rect 89374 550170 89442 550226
rect 89498 550170 120038 550226
rect 120094 550170 120162 550226
rect 120218 550170 150758 550226
rect 150814 550170 150882 550226
rect 150938 550170 181478 550226
rect 181534 550170 181602 550226
rect 181658 550170 212198 550226
rect 212254 550170 212322 550226
rect 212378 550170 242918 550226
rect 242974 550170 243042 550226
rect 243098 550170 273638 550226
rect 273694 550170 273762 550226
rect 273818 550170 304358 550226
rect 304414 550170 304482 550226
rect 304538 550170 335078 550226
rect 335134 550170 335202 550226
rect 335258 550170 365798 550226
rect 365854 550170 365922 550226
rect 365978 550170 396518 550226
rect 396574 550170 396642 550226
rect 396698 550170 427238 550226
rect 427294 550170 427362 550226
rect 427418 550170 457958 550226
rect 458014 550170 458082 550226
rect 458138 550170 488678 550226
rect 488734 550170 488802 550226
rect 488858 550170 519398 550226
rect 519454 550170 519522 550226
rect 519578 550170 550118 550226
rect 550174 550170 550242 550226
rect 550298 550170 592914 550226
rect 592970 550170 593038 550226
rect 593094 550170 593162 550226
rect 593218 550170 593286 550226
rect 593342 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect -1916 550102 597980 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 27878 550102
rect 27934 550046 28002 550102
rect 28058 550046 58598 550102
rect 58654 550046 58722 550102
rect 58778 550046 89318 550102
rect 89374 550046 89442 550102
rect 89498 550046 120038 550102
rect 120094 550046 120162 550102
rect 120218 550046 150758 550102
rect 150814 550046 150882 550102
rect 150938 550046 181478 550102
rect 181534 550046 181602 550102
rect 181658 550046 212198 550102
rect 212254 550046 212322 550102
rect 212378 550046 242918 550102
rect 242974 550046 243042 550102
rect 243098 550046 273638 550102
rect 273694 550046 273762 550102
rect 273818 550046 304358 550102
rect 304414 550046 304482 550102
rect 304538 550046 335078 550102
rect 335134 550046 335202 550102
rect 335258 550046 365798 550102
rect 365854 550046 365922 550102
rect 365978 550046 396518 550102
rect 396574 550046 396642 550102
rect 396698 550046 427238 550102
rect 427294 550046 427362 550102
rect 427418 550046 457958 550102
rect 458014 550046 458082 550102
rect 458138 550046 488678 550102
rect 488734 550046 488802 550102
rect 488858 550046 519398 550102
rect 519454 550046 519522 550102
rect 519578 550046 550118 550102
rect 550174 550046 550242 550102
rect 550298 550046 592914 550102
rect 592970 550046 593038 550102
rect 593094 550046 593162 550102
rect 593218 550046 593286 550102
rect 593342 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect -1916 549978 597980 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 27878 549978
rect 27934 549922 28002 549978
rect 28058 549922 58598 549978
rect 58654 549922 58722 549978
rect 58778 549922 89318 549978
rect 89374 549922 89442 549978
rect 89498 549922 120038 549978
rect 120094 549922 120162 549978
rect 120218 549922 150758 549978
rect 150814 549922 150882 549978
rect 150938 549922 181478 549978
rect 181534 549922 181602 549978
rect 181658 549922 212198 549978
rect 212254 549922 212322 549978
rect 212378 549922 242918 549978
rect 242974 549922 243042 549978
rect 243098 549922 273638 549978
rect 273694 549922 273762 549978
rect 273818 549922 304358 549978
rect 304414 549922 304482 549978
rect 304538 549922 335078 549978
rect 335134 549922 335202 549978
rect 335258 549922 365798 549978
rect 365854 549922 365922 549978
rect 365978 549922 396518 549978
rect 396574 549922 396642 549978
rect 396698 549922 427238 549978
rect 427294 549922 427362 549978
rect 427418 549922 457958 549978
rect 458014 549922 458082 549978
rect 458138 549922 488678 549978
rect 488734 549922 488802 549978
rect 488858 549922 519398 549978
rect 519454 549922 519522 549978
rect 519578 549922 550118 549978
rect 550174 549922 550242 549978
rect 550298 549922 592914 549978
rect 592970 549922 593038 549978
rect 593094 549922 593162 549978
rect 593218 549922 593286 549978
rect 593342 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect -1916 549826 597980 549922
rect -1916 544350 597980 544446
rect -1916 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 5514 544350
rect 5570 544294 5638 544350
rect 5694 544294 5762 544350
rect 5818 544294 5886 544350
rect 5942 544294 12518 544350
rect 12574 544294 12642 544350
rect 12698 544294 43238 544350
rect 43294 544294 43362 544350
rect 43418 544294 73958 544350
rect 74014 544294 74082 544350
rect 74138 544294 104678 544350
rect 104734 544294 104802 544350
rect 104858 544294 135398 544350
rect 135454 544294 135522 544350
rect 135578 544294 166118 544350
rect 166174 544294 166242 544350
rect 166298 544294 196838 544350
rect 196894 544294 196962 544350
rect 197018 544294 227558 544350
rect 227614 544294 227682 544350
rect 227738 544294 258278 544350
rect 258334 544294 258402 544350
rect 258458 544294 288998 544350
rect 289054 544294 289122 544350
rect 289178 544294 319718 544350
rect 319774 544294 319842 544350
rect 319898 544294 350438 544350
rect 350494 544294 350562 544350
rect 350618 544294 381158 544350
rect 381214 544294 381282 544350
rect 381338 544294 411878 544350
rect 411934 544294 412002 544350
rect 412058 544294 442598 544350
rect 442654 544294 442722 544350
rect 442778 544294 473318 544350
rect 473374 544294 473442 544350
rect 473498 544294 504038 544350
rect 504094 544294 504162 544350
rect 504218 544294 534758 544350
rect 534814 544294 534882 544350
rect 534938 544294 565478 544350
rect 565534 544294 565602 544350
rect 565658 544294 589194 544350
rect 589250 544294 589318 544350
rect 589374 544294 589442 544350
rect 589498 544294 589566 544350
rect 589622 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597980 544350
rect -1916 544226 597980 544294
rect -1916 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 5514 544226
rect 5570 544170 5638 544226
rect 5694 544170 5762 544226
rect 5818 544170 5886 544226
rect 5942 544170 12518 544226
rect 12574 544170 12642 544226
rect 12698 544170 43238 544226
rect 43294 544170 43362 544226
rect 43418 544170 73958 544226
rect 74014 544170 74082 544226
rect 74138 544170 104678 544226
rect 104734 544170 104802 544226
rect 104858 544170 135398 544226
rect 135454 544170 135522 544226
rect 135578 544170 166118 544226
rect 166174 544170 166242 544226
rect 166298 544170 196838 544226
rect 196894 544170 196962 544226
rect 197018 544170 227558 544226
rect 227614 544170 227682 544226
rect 227738 544170 258278 544226
rect 258334 544170 258402 544226
rect 258458 544170 288998 544226
rect 289054 544170 289122 544226
rect 289178 544170 319718 544226
rect 319774 544170 319842 544226
rect 319898 544170 350438 544226
rect 350494 544170 350562 544226
rect 350618 544170 381158 544226
rect 381214 544170 381282 544226
rect 381338 544170 411878 544226
rect 411934 544170 412002 544226
rect 412058 544170 442598 544226
rect 442654 544170 442722 544226
rect 442778 544170 473318 544226
rect 473374 544170 473442 544226
rect 473498 544170 504038 544226
rect 504094 544170 504162 544226
rect 504218 544170 534758 544226
rect 534814 544170 534882 544226
rect 534938 544170 565478 544226
rect 565534 544170 565602 544226
rect 565658 544170 589194 544226
rect 589250 544170 589318 544226
rect 589374 544170 589442 544226
rect 589498 544170 589566 544226
rect 589622 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597980 544226
rect -1916 544102 597980 544170
rect -1916 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 5514 544102
rect 5570 544046 5638 544102
rect 5694 544046 5762 544102
rect 5818 544046 5886 544102
rect 5942 544046 12518 544102
rect 12574 544046 12642 544102
rect 12698 544046 43238 544102
rect 43294 544046 43362 544102
rect 43418 544046 73958 544102
rect 74014 544046 74082 544102
rect 74138 544046 104678 544102
rect 104734 544046 104802 544102
rect 104858 544046 135398 544102
rect 135454 544046 135522 544102
rect 135578 544046 166118 544102
rect 166174 544046 166242 544102
rect 166298 544046 196838 544102
rect 196894 544046 196962 544102
rect 197018 544046 227558 544102
rect 227614 544046 227682 544102
rect 227738 544046 258278 544102
rect 258334 544046 258402 544102
rect 258458 544046 288998 544102
rect 289054 544046 289122 544102
rect 289178 544046 319718 544102
rect 319774 544046 319842 544102
rect 319898 544046 350438 544102
rect 350494 544046 350562 544102
rect 350618 544046 381158 544102
rect 381214 544046 381282 544102
rect 381338 544046 411878 544102
rect 411934 544046 412002 544102
rect 412058 544046 442598 544102
rect 442654 544046 442722 544102
rect 442778 544046 473318 544102
rect 473374 544046 473442 544102
rect 473498 544046 504038 544102
rect 504094 544046 504162 544102
rect 504218 544046 534758 544102
rect 534814 544046 534882 544102
rect 534938 544046 565478 544102
rect 565534 544046 565602 544102
rect 565658 544046 589194 544102
rect 589250 544046 589318 544102
rect 589374 544046 589442 544102
rect 589498 544046 589566 544102
rect 589622 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597980 544102
rect -1916 543978 597980 544046
rect -1916 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 5514 543978
rect 5570 543922 5638 543978
rect 5694 543922 5762 543978
rect 5818 543922 5886 543978
rect 5942 543922 12518 543978
rect 12574 543922 12642 543978
rect 12698 543922 43238 543978
rect 43294 543922 43362 543978
rect 43418 543922 73958 543978
rect 74014 543922 74082 543978
rect 74138 543922 104678 543978
rect 104734 543922 104802 543978
rect 104858 543922 135398 543978
rect 135454 543922 135522 543978
rect 135578 543922 166118 543978
rect 166174 543922 166242 543978
rect 166298 543922 196838 543978
rect 196894 543922 196962 543978
rect 197018 543922 227558 543978
rect 227614 543922 227682 543978
rect 227738 543922 258278 543978
rect 258334 543922 258402 543978
rect 258458 543922 288998 543978
rect 289054 543922 289122 543978
rect 289178 543922 319718 543978
rect 319774 543922 319842 543978
rect 319898 543922 350438 543978
rect 350494 543922 350562 543978
rect 350618 543922 381158 543978
rect 381214 543922 381282 543978
rect 381338 543922 411878 543978
rect 411934 543922 412002 543978
rect 412058 543922 442598 543978
rect 442654 543922 442722 543978
rect 442778 543922 473318 543978
rect 473374 543922 473442 543978
rect 473498 543922 504038 543978
rect 504094 543922 504162 543978
rect 504218 543922 534758 543978
rect 534814 543922 534882 543978
rect 534938 543922 565478 543978
rect 565534 543922 565602 543978
rect 565658 543922 589194 543978
rect 589250 543922 589318 543978
rect 589374 543922 589442 543978
rect 589498 543922 589566 543978
rect 589622 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597980 543978
rect -1916 543826 597980 543922
rect -1916 532350 597980 532446
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 27878 532350
rect 27934 532294 28002 532350
rect 28058 532294 58598 532350
rect 58654 532294 58722 532350
rect 58778 532294 89318 532350
rect 89374 532294 89442 532350
rect 89498 532294 120038 532350
rect 120094 532294 120162 532350
rect 120218 532294 150758 532350
rect 150814 532294 150882 532350
rect 150938 532294 181478 532350
rect 181534 532294 181602 532350
rect 181658 532294 212198 532350
rect 212254 532294 212322 532350
rect 212378 532294 242918 532350
rect 242974 532294 243042 532350
rect 243098 532294 273638 532350
rect 273694 532294 273762 532350
rect 273818 532294 304358 532350
rect 304414 532294 304482 532350
rect 304538 532294 335078 532350
rect 335134 532294 335202 532350
rect 335258 532294 365798 532350
rect 365854 532294 365922 532350
rect 365978 532294 396518 532350
rect 396574 532294 396642 532350
rect 396698 532294 427238 532350
rect 427294 532294 427362 532350
rect 427418 532294 457958 532350
rect 458014 532294 458082 532350
rect 458138 532294 488678 532350
rect 488734 532294 488802 532350
rect 488858 532294 519398 532350
rect 519454 532294 519522 532350
rect 519578 532294 550118 532350
rect 550174 532294 550242 532350
rect 550298 532294 592914 532350
rect 592970 532294 593038 532350
rect 593094 532294 593162 532350
rect 593218 532294 593286 532350
rect 593342 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect -1916 532226 597980 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 27878 532226
rect 27934 532170 28002 532226
rect 28058 532170 58598 532226
rect 58654 532170 58722 532226
rect 58778 532170 89318 532226
rect 89374 532170 89442 532226
rect 89498 532170 120038 532226
rect 120094 532170 120162 532226
rect 120218 532170 150758 532226
rect 150814 532170 150882 532226
rect 150938 532170 181478 532226
rect 181534 532170 181602 532226
rect 181658 532170 212198 532226
rect 212254 532170 212322 532226
rect 212378 532170 242918 532226
rect 242974 532170 243042 532226
rect 243098 532170 273638 532226
rect 273694 532170 273762 532226
rect 273818 532170 304358 532226
rect 304414 532170 304482 532226
rect 304538 532170 335078 532226
rect 335134 532170 335202 532226
rect 335258 532170 365798 532226
rect 365854 532170 365922 532226
rect 365978 532170 396518 532226
rect 396574 532170 396642 532226
rect 396698 532170 427238 532226
rect 427294 532170 427362 532226
rect 427418 532170 457958 532226
rect 458014 532170 458082 532226
rect 458138 532170 488678 532226
rect 488734 532170 488802 532226
rect 488858 532170 519398 532226
rect 519454 532170 519522 532226
rect 519578 532170 550118 532226
rect 550174 532170 550242 532226
rect 550298 532170 592914 532226
rect 592970 532170 593038 532226
rect 593094 532170 593162 532226
rect 593218 532170 593286 532226
rect 593342 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect -1916 532102 597980 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 27878 532102
rect 27934 532046 28002 532102
rect 28058 532046 58598 532102
rect 58654 532046 58722 532102
rect 58778 532046 89318 532102
rect 89374 532046 89442 532102
rect 89498 532046 120038 532102
rect 120094 532046 120162 532102
rect 120218 532046 150758 532102
rect 150814 532046 150882 532102
rect 150938 532046 181478 532102
rect 181534 532046 181602 532102
rect 181658 532046 212198 532102
rect 212254 532046 212322 532102
rect 212378 532046 242918 532102
rect 242974 532046 243042 532102
rect 243098 532046 273638 532102
rect 273694 532046 273762 532102
rect 273818 532046 304358 532102
rect 304414 532046 304482 532102
rect 304538 532046 335078 532102
rect 335134 532046 335202 532102
rect 335258 532046 365798 532102
rect 365854 532046 365922 532102
rect 365978 532046 396518 532102
rect 396574 532046 396642 532102
rect 396698 532046 427238 532102
rect 427294 532046 427362 532102
rect 427418 532046 457958 532102
rect 458014 532046 458082 532102
rect 458138 532046 488678 532102
rect 488734 532046 488802 532102
rect 488858 532046 519398 532102
rect 519454 532046 519522 532102
rect 519578 532046 550118 532102
rect 550174 532046 550242 532102
rect 550298 532046 592914 532102
rect 592970 532046 593038 532102
rect 593094 532046 593162 532102
rect 593218 532046 593286 532102
rect 593342 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect -1916 531978 597980 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 27878 531978
rect 27934 531922 28002 531978
rect 28058 531922 58598 531978
rect 58654 531922 58722 531978
rect 58778 531922 89318 531978
rect 89374 531922 89442 531978
rect 89498 531922 120038 531978
rect 120094 531922 120162 531978
rect 120218 531922 150758 531978
rect 150814 531922 150882 531978
rect 150938 531922 181478 531978
rect 181534 531922 181602 531978
rect 181658 531922 212198 531978
rect 212254 531922 212322 531978
rect 212378 531922 242918 531978
rect 242974 531922 243042 531978
rect 243098 531922 273638 531978
rect 273694 531922 273762 531978
rect 273818 531922 304358 531978
rect 304414 531922 304482 531978
rect 304538 531922 335078 531978
rect 335134 531922 335202 531978
rect 335258 531922 365798 531978
rect 365854 531922 365922 531978
rect 365978 531922 396518 531978
rect 396574 531922 396642 531978
rect 396698 531922 427238 531978
rect 427294 531922 427362 531978
rect 427418 531922 457958 531978
rect 458014 531922 458082 531978
rect 458138 531922 488678 531978
rect 488734 531922 488802 531978
rect 488858 531922 519398 531978
rect 519454 531922 519522 531978
rect 519578 531922 550118 531978
rect 550174 531922 550242 531978
rect 550298 531922 592914 531978
rect 592970 531922 593038 531978
rect 593094 531922 593162 531978
rect 593218 531922 593286 531978
rect 593342 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect -1916 531826 597980 531922
rect -1916 526350 597980 526446
rect -1916 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 5514 526350
rect 5570 526294 5638 526350
rect 5694 526294 5762 526350
rect 5818 526294 5886 526350
rect 5942 526294 12518 526350
rect 12574 526294 12642 526350
rect 12698 526294 43238 526350
rect 43294 526294 43362 526350
rect 43418 526294 73958 526350
rect 74014 526294 74082 526350
rect 74138 526294 104678 526350
rect 104734 526294 104802 526350
rect 104858 526294 135398 526350
rect 135454 526294 135522 526350
rect 135578 526294 166118 526350
rect 166174 526294 166242 526350
rect 166298 526294 196838 526350
rect 196894 526294 196962 526350
rect 197018 526294 227558 526350
rect 227614 526294 227682 526350
rect 227738 526294 258278 526350
rect 258334 526294 258402 526350
rect 258458 526294 288998 526350
rect 289054 526294 289122 526350
rect 289178 526294 319718 526350
rect 319774 526294 319842 526350
rect 319898 526294 350438 526350
rect 350494 526294 350562 526350
rect 350618 526294 381158 526350
rect 381214 526294 381282 526350
rect 381338 526294 411878 526350
rect 411934 526294 412002 526350
rect 412058 526294 442598 526350
rect 442654 526294 442722 526350
rect 442778 526294 473318 526350
rect 473374 526294 473442 526350
rect 473498 526294 504038 526350
rect 504094 526294 504162 526350
rect 504218 526294 534758 526350
rect 534814 526294 534882 526350
rect 534938 526294 565478 526350
rect 565534 526294 565602 526350
rect 565658 526294 589194 526350
rect 589250 526294 589318 526350
rect 589374 526294 589442 526350
rect 589498 526294 589566 526350
rect 589622 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597980 526350
rect -1916 526226 597980 526294
rect -1916 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 5514 526226
rect 5570 526170 5638 526226
rect 5694 526170 5762 526226
rect 5818 526170 5886 526226
rect 5942 526170 12518 526226
rect 12574 526170 12642 526226
rect 12698 526170 43238 526226
rect 43294 526170 43362 526226
rect 43418 526170 73958 526226
rect 74014 526170 74082 526226
rect 74138 526170 104678 526226
rect 104734 526170 104802 526226
rect 104858 526170 135398 526226
rect 135454 526170 135522 526226
rect 135578 526170 166118 526226
rect 166174 526170 166242 526226
rect 166298 526170 196838 526226
rect 196894 526170 196962 526226
rect 197018 526170 227558 526226
rect 227614 526170 227682 526226
rect 227738 526170 258278 526226
rect 258334 526170 258402 526226
rect 258458 526170 288998 526226
rect 289054 526170 289122 526226
rect 289178 526170 319718 526226
rect 319774 526170 319842 526226
rect 319898 526170 350438 526226
rect 350494 526170 350562 526226
rect 350618 526170 381158 526226
rect 381214 526170 381282 526226
rect 381338 526170 411878 526226
rect 411934 526170 412002 526226
rect 412058 526170 442598 526226
rect 442654 526170 442722 526226
rect 442778 526170 473318 526226
rect 473374 526170 473442 526226
rect 473498 526170 504038 526226
rect 504094 526170 504162 526226
rect 504218 526170 534758 526226
rect 534814 526170 534882 526226
rect 534938 526170 565478 526226
rect 565534 526170 565602 526226
rect 565658 526170 589194 526226
rect 589250 526170 589318 526226
rect 589374 526170 589442 526226
rect 589498 526170 589566 526226
rect 589622 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597980 526226
rect -1916 526102 597980 526170
rect -1916 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 5514 526102
rect 5570 526046 5638 526102
rect 5694 526046 5762 526102
rect 5818 526046 5886 526102
rect 5942 526046 12518 526102
rect 12574 526046 12642 526102
rect 12698 526046 43238 526102
rect 43294 526046 43362 526102
rect 43418 526046 73958 526102
rect 74014 526046 74082 526102
rect 74138 526046 104678 526102
rect 104734 526046 104802 526102
rect 104858 526046 135398 526102
rect 135454 526046 135522 526102
rect 135578 526046 166118 526102
rect 166174 526046 166242 526102
rect 166298 526046 196838 526102
rect 196894 526046 196962 526102
rect 197018 526046 227558 526102
rect 227614 526046 227682 526102
rect 227738 526046 258278 526102
rect 258334 526046 258402 526102
rect 258458 526046 288998 526102
rect 289054 526046 289122 526102
rect 289178 526046 319718 526102
rect 319774 526046 319842 526102
rect 319898 526046 350438 526102
rect 350494 526046 350562 526102
rect 350618 526046 381158 526102
rect 381214 526046 381282 526102
rect 381338 526046 411878 526102
rect 411934 526046 412002 526102
rect 412058 526046 442598 526102
rect 442654 526046 442722 526102
rect 442778 526046 473318 526102
rect 473374 526046 473442 526102
rect 473498 526046 504038 526102
rect 504094 526046 504162 526102
rect 504218 526046 534758 526102
rect 534814 526046 534882 526102
rect 534938 526046 565478 526102
rect 565534 526046 565602 526102
rect 565658 526046 589194 526102
rect 589250 526046 589318 526102
rect 589374 526046 589442 526102
rect 589498 526046 589566 526102
rect 589622 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597980 526102
rect -1916 525978 597980 526046
rect -1916 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 5514 525978
rect 5570 525922 5638 525978
rect 5694 525922 5762 525978
rect 5818 525922 5886 525978
rect 5942 525922 12518 525978
rect 12574 525922 12642 525978
rect 12698 525922 43238 525978
rect 43294 525922 43362 525978
rect 43418 525922 73958 525978
rect 74014 525922 74082 525978
rect 74138 525922 104678 525978
rect 104734 525922 104802 525978
rect 104858 525922 135398 525978
rect 135454 525922 135522 525978
rect 135578 525922 166118 525978
rect 166174 525922 166242 525978
rect 166298 525922 196838 525978
rect 196894 525922 196962 525978
rect 197018 525922 227558 525978
rect 227614 525922 227682 525978
rect 227738 525922 258278 525978
rect 258334 525922 258402 525978
rect 258458 525922 288998 525978
rect 289054 525922 289122 525978
rect 289178 525922 319718 525978
rect 319774 525922 319842 525978
rect 319898 525922 350438 525978
rect 350494 525922 350562 525978
rect 350618 525922 381158 525978
rect 381214 525922 381282 525978
rect 381338 525922 411878 525978
rect 411934 525922 412002 525978
rect 412058 525922 442598 525978
rect 442654 525922 442722 525978
rect 442778 525922 473318 525978
rect 473374 525922 473442 525978
rect 473498 525922 504038 525978
rect 504094 525922 504162 525978
rect 504218 525922 534758 525978
rect 534814 525922 534882 525978
rect 534938 525922 565478 525978
rect 565534 525922 565602 525978
rect 565658 525922 589194 525978
rect 589250 525922 589318 525978
rect 589374 525922 589442 525978
rect 589498 525922 589566 525978
rect 589622 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597980 525978
rect -1916 525826 597980 525922
rect -1916 514350 597980 514446
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 27878 514350
rect 27934 514294 28002 514350
rect 28058 514294 58598 514350
rect 58654 514294 58722 514350
rect 58778 514294 89318 514350
rect 89374 514294 89442 514350
rect 89498 514294 120038 514350
rect 120094 514294 120162 514350
rect 120218 514294 150758 514350
rect 150814 514294 150882 514350
rect 150938 514294 181478 514350
rect 181534 514294 181602 514350
rect 181658 514294 212198 514350
rect 212254 514294 212322 514350
rect 212378 514294 242918 514350
rect 242974 514294 243042 514350
rect 243098 514294 273638 514350
rect 273694 514294 273762 514350
rect 273818 514294 304358 514350
rect 304414 514294 304482 514350
rect 304538 514294 335078 514350
rect 335134 514294 335202 514350
rect 335258 514294 365798 514350
rect 365854 514294 365922 514350
rect 365978 514294 396518 514350
rect 396574 514294 396642 514350
rect 396698 514294 427238 514350
rect 427294 514294 427362 514350
rect 427418 514294 457958 514350
rect 458014 514294 458082 514350
rect 458138 514294 488678 514350
rect 488734 514294 488802 514350
rect 488858 514294 519398 514350
rect 519454 514294 519522 514350
rect 519578 514294 550118 514350
rect 550174 514294 550242 514350
rect 550298 514294 592914 514350
rect 592970 514294 593038 514350
rect 593094 514294 593162 514350
rect 593218 514294 593286 514350
rect 593342 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect -1916 514226 597980 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 27878 514226
rect 27934 514170 28002 514226
rect 28058 514170 58598 514226
rect 58654 514170 58722 514226
rect 58778 514170 89318 514226
rect 89374 514170 89442 514226
rect 89498 514170 120038 514226
rect 120094 514170 120162 514226
rect 120218 514170 150758 514226
rect 150814 514170 150882 514226
rect 150938 514170 181478 514226
rect 181534 514170 181602 514226
rect 181658 514170 212198 514226
rect 212254 514170 212322 514226
rect 212378 514170 242918 514226
rect 242974 514170 243042 514226
rect 243098 514170 273638 514226
rect 273694 514170 273762 514226
rect 273818 514170 304358 514226
rect 304414 514170 304482 514226
rect 304538 514170 335078 514226
rect 335134 514170 335202 514226
rect 335258 514170 365798 514226
rect 365854 514170 365922 514226
rect 365978 514170 396518 514226
rect 396574 514170 396642 514226
rect 396698 514170 427238 514226
rect 427294 514170 427362 514226
rect 427418 514170 457958 514226
rect 458014 514170 458082 514226
rect 458138 514170 488678 514226
rect 488734 514170 488802 514226
rect 488858 514170 519398 514226
rect 519454 514170 519522 514226
rect 519578 514170 550118 514226
rect 550174 514170 550242 514226
rect 550298 514170 592914 514226
rect 592970 514170 593038 514226
rect 593094 514170 593162 514226
rect 593218 514170 593286 514226
rect 593342 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect -1916 514102 597980 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 27878 514102
rect 27934 514046 28002 514102
rect 28058 514046 58598 514102
rect 58654 514046 58722 514102
rect 58778 514046 89318 514102
rect 89374 514046 89442 514102
rect 89498 514046 120038 514102
rect 120094 514046 120162 514102
rect 120218 514046 150758 514102
rect 150814 514046 150882 514102
rect 150938 514046 181478 514102
rect 181534 514046 181602 514102
rect 181658 514046 212198 514102
rect 212254 514046 212322 514102
rect 212378 514046 242918 514102
rect 242974 514046 243042 514102
rect 243098 514046 273638 514102
rect 273694 514046 273762 514102
rect 273818 514046 304358 514102
rect 304414 514046 304482 514102
rect 304538 514046 335078 514102
rect 335134 514046 335202 514102
rect 335258 514046 365798 514102
rect 365854 514046 365922 514102
rect 365978 514046 396518 514102
rect 396574 514046 396642 514102
rect 396698 514046 427238 514102
rect 427294 514046 427362 514102
rect 427418 514046 457958 514102
rect 458014 514046 458082 514102
rect 458138 514046 488678 514102
rect 488734 514046 488802 514102
rect 488858 514046 519398 514102
rect 519454 514046 519522 514102
rect 519578 514046 550118 514102
rect 550174 514046 550242 514102
rect 550298 514046 592914 514102
rect 592970 514046 593038 514102
rect 593094 514046 593162 514102
rect 593218 514046 593286 514102
rect 593342 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect -1916 513978 597980 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 27878 513978
rect 27934 513922 28002 513978
rect 28058 513922 58598 513978
rect 58654 513922 58722 513978
rect 58778 513922 89318 513978
rect 89374 513922 89442 513978
rect 89498 513922 120038 513978
rect 120094 513922 120162 513978
rect 120218 513922 150758 513978
rect 150814 513922 150882 513978
rect 150938 513922 181478 513978
rect 181534 513922 181602 513978
rect 181658 513922 212198 513978
rect 212254 513922 212322 513978
rect 212378 513922 242918 513978
rect 242974 513922 243042 513978
rect 243098 513922 273638 513978
rect 273694 513922 273762 513978
rect 273818 513922 304358 513978
rect 304414 513922 304482 513978
rect 304538 513922 335078 513978
rect 335134 513922 335202 513978
rect 335258 513922 365798 513978
rect 365854 513922 365922 513978
rect 365978 513922 396518 513978
rect 396574 513922 396642 513978
rect 396698 513922 427238 513978
rect 427294 513922 427362 513978
rect 427418 513922 457958 513978
rect 458014 513922 458082 513978
rect 458138 513922 488678 513978
rect 488734 513922 488802 513978
rect 488858 513922 519398 513978
rect 519454 513922 519522 513978
rect 519578 513922 550118 513978
rect 550174 513922 550242 513978
rect 550298 513922 592914 513978
rect 592970 513922 593038 513978
rect 593094 513922 593162 513978
rect 593218 513922 593286 513978
rect 593342 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect -1916 513826 597980 513922
rect -1916 508350 597980 508446
rect -1916 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 5514 508350
rect 5570 508294 5638 508350
rect 5694 508294 5762 508350
rect 5818 508294 5886 508350
rect 5942 508294 12518 508350
rect 12574 508294 12642 508350
rect 12698 508294 43238 508350
rect 43294 508294 43362 508350
rect 43418 508294 73958 508350
rect 74014 508294 74082 508350
rect 74138 508294 104678 508350
rect 104734 508294 104802 508350
rect 104858 508294 135398 508350
rect 135454 508294 135522 508350
rect 135578 508294 166118 508350
rect 166174 508294 166242 508350
rect 166298 508294 196838 508350
rect 196894 508294 196962 508350
rect 197018 508294 227558 508350
rect 227614 508294 227682 508350
rect 227738 508294 258278 508350
rect 258334 508294 258402 508350
rect 258458 508294 288998 508350
rect 289054 508294 289122 508350
rect 289178 508294 319718 508350
rect 319774 508294 319842 508350
rect 319898 508294 350438 508350
rect 350494 508294 350562 508350
rect 350618 508294 381158 508350
rect 381214 508294 381282 508350
rect 381338 508294 411878 508350
rect 411934 508294 412002 508350
rect 412058 508294 442598 508350
rect 442654 508294 442722 508350
rect 442778 508294 473318 508350
rect 473374 508294 473442 508350
rect 473498 508294 504038 508350
rect 504094 508294 504162 508350
rect 504218 508294 534758 508350
rect 534814 508294 534882 508350
rect 534938 508294 565478 508350
rect 565534 508294 565602 508350
rect 565658 508294 589194 508350
rect 589250 508294 589318 508350
rect 589374 508294 589442 508350
rect 589498 508294 589566 508350
rect 589622 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597980 508350
rect -1916 508226 597980 508294
rect -1916 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 5514 508226
rect 5570 508170 5638 508226
rect 5694 508170 5762 508226
rect 5818 508170 5886 508226
rect 5942 508170 12518 508226
rect 12574 508170 12642 508226
rect 12698 508170 43238 508226
rect 43294 508170 43362 508226
rect 43418 508170 73958 508226
rect 74014 508170 74082 508226
rect 74138 508170 104678 508226
rect 104734 508170 104802 508226
rect 104858 508170 135398 508226
rect 135454 508170 135522 508226
rect 135578 508170 166118 508226
rect 166174 508170 166242 508226
rect 166298 508170 196838 508226
rect 196894 508170 196962 508226
rect 197018 508170 227558 508226
rect 227614 508170 227682 508226
rect 227738 508170 258278 508226
rect 258334 508170 258402 508226
rect 258458 508170 288998 508226
rect 289054 508170 289122 508226
rect 289178 508170 319718 508226
rect 319774 508170 319842 508226
rect 319898 508170 350438 508226
rect 350494 508170 350562 508226
rect 350618 508170 381158 508226
rect 381214 508170 381282 508226
rect 381338 508170 411878 508226
rect 411934 508170 412002 508226
rect 412058 508170 442598 508226
rect 442654 508170 442722 508226
rect 442778 508170 473318 508226
rect 473374 508170 473442 508226
rect 473498 508170 504038 508226
rect 504094 508170 504162 508226
rect 504218 508170 534758 508226
rect 534814 508170 534882 508226
rect 534938 508170 565478 508226
rect 565534 508170 565602 508226
rect 565658 508170 589194 508226
rect 589250 508170 589318 508226
rect 589374 508170 589442 508226
rect 589498 508170 589566 508226
rect 589622 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597980 508226
rect -1916 508102 597980 508170
rect -1916 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 5514 508102
rect 5570 508046 5638 508102
rect 5694 508046 5762 508102
rect 5818 508046 5886 508102
rect 5942 508046 12518 508102
rect 12574 508046 12642 508102
rect 12698 508046 43238 508102
rect 43294 508046 43362 508102
rect 43418 508046 73958 508102
rect 74014 508046 74082 508102
rect 74138 508046 104678 508102
rect 104734 508046 104802 508102
rect 104858 508046 135398 508102
rect 135454 508046 135522 508102
rect 135578 508046 166118 508102
rect 166174 508046 166242 508102
rect 166298 508046 196838 508102
rect 196894 508046 196962 508102
rect 197018 508046 227558 508102
rect 227614 508046 227682 508102
rect 227738 508046 258278 508102
rect 258334 508046 258402 508102
rect 258458 508046 288998 508102
rect 289054 508046 289122 508102
rect 289178 508046 319718 508102
rect 319774 508046 319842 508102
rect 319898 508046 350438 508102
rect 350494 508046 350562 508102
rect 350618 508046 381158 508102
rect 381214 508046 381282 508102
rect 381338 508046 411878 508102
rect 411934 508046 412002 508102
rect 412058 508046 442598 508102
rect 442654 508046 442722 508102
rect 442778 508046 473318 508102
rect 473374 508046 473442 508102
rect 473498 508046 504038 508102
rect 504094 508046 504162 508102
rect 504218 508046 534758 508102
rect 534814 508046 534882 508102
rect 534938 508046 565478 508102
rect 565534 508046 565602 508102
rect 565658 508046 589194 508102
rect 589250 508046 589318 508102
rect 589374 508046 589442 508102
rect 589498 508046 589566 508102
rect 589622 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597980 508102
rect -1916 507978 597980 508046
rect -1916 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 5514 507978
rect 5570 507922 5638 507978
rect 5694 507922 5762 507978
rect 5818 507922 5886 507978
rect 5942 507922 12518 507978
rect 12574 507922 12642 507978
rect 12698 507922 43238 507978
rect 43294 507922 43362 507978
rect 43418 507922 73958 507978
rect 74014 507922 74082 507978
rect 74138 507922 104678 507978
rect 104734 507922 104802 507978
rect 104858 507922 135398 507978
rect 135454 507922 135522 507978
rect 135578 507922 166118 507978
rect 166174 507922 166242 507978
rect 166298 507922 196838 507978
rect 196894 507922 196962 507978
rect 197018 507922 227558 507978
rect 227614 507922 227682 507978
rect 227738 507922 258278 507978
rect 258334 507922 258402 507978
rect 258458 507922 288998 507978
rect 289054 507922 289122 507978
rect 289178 507922 319718 507978
rect 319774 507922 319842 507978
rect 319898 507922 350438 507978
rect 350494 507922 350562 507978
rect 350618 507922 381158 507978
rect 381214 507922 381282 507978
rect 381338 507922 411878 507978
rect 411934 507922 412002 507978
rect 412058 507922 442598 507978
rect 442654 507922 442722 507978
rect 442778 507922 473318 507978
rect 473374 507922 473442 507978
rect 473498 507922 504038 507978
rect 504094 507922 504162 507978
rect 504218 507922 534758 507978
rect 534814 507922 534882 507978
rect 534938 507922 565478 507978
rect 565534 507922 565602 507978
rect 565658 507922 589194 507978
rect 589250 507922 589318 507978
rect 589374 507922 589442 507978
rect 589498 507922 589566 507978
rect 589622 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597980 507978
rect -1916 507826 597980 507922
rect -1916 496350 597980 496446
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 27878 496350
rect 27934 496294 28002 496350
rect 28058 496294 58598 496350
rect 58654 496294 58722 496350
rect 58778 496294 89318 496350
rect 89374 496294 89442 496350
rect 89498 496294 120038 496350
rect 120094 496294 120162 496350
rect 120218 496294 150758 496350
rect 150814 496294 150882 496350
rect 150938 496294 181478 496350
rect 181534 496294 181602 496350
rect 181658 496294 212198 496350
rect 212254 496294 212322 496350
rect 212378 496294 242918 496350
rect 242974 496294 243042 496350
rect 243098 496294 273638 496350
rect 273694 496294 273762 496350
rect 273818 496294 304358 496350
rect 304414 496294 304482 496350
rect 304538 496294 335078 496350
rect 335134 496294 335202 496350
rect 335258 496294 365798 496350
rect 365854 496294 365922 496350
rect 365978 496294 396518 496350
rect 396574 496294 396642 496350
rect 396698 496294 427238 496350
rect 427294 496294 427362 496350
rect 427418 496294 457958 496350
rect 458014 496294 458082 496350
rect 458138 496294 488678 496350
rect 488734 496294 488802 496350
rect 488858 496294 519398 496350
rect 519454 496294 519522 496350
rect 519578 496294 550118 496350
rect 550174 496294 550242 496350
rect 550298 496294 592914 496350
rect 592970 496294 593038 496350
rect 593094 496294 593162 496350
rect 593218 496294 593286 496350
rect 593342 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect -1916 496226 597980 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 27878 496226
rect 27934 496170 28002 496226
rect 28058 496170 58598 496226
rect 58654 496170 58722 496226
rect 58778 496170 89318 496226
rect 89374 496170 89442 496226
rect 89498 496170 120038 496226
rect 120094 496170 120162 496226
rect 120218 496170 150758 496226
rect 150814 496170 150882 496226
rect 150938 496170 181478 496226
rect 181534 496170 181602 496226
rect 181658 496170 212198 496226
rect 212254 496170 212322 496226
rect 212378 496170 242918 496226
rect 242974 496170 243042 496226
rect 243098 496170 273638 496226
rect 273694 496170 273762 496226
rect 273818 496170 304358 496226
rect 304414 496170 304482 496226
rect 304538 496170 335078 496226
rect 335134 496170 335202 496226
rect 335258 496170 365798 496226
rect 365854 496170 365922 496226
rect 365978 496170 396518 496226
rect 396574 496170 396642 496226
rect 396698 496170 427238 496226
rect 427294 496170 427362 496226
rect 427418 496170 457958 496226
rect 458014 496170 458082 496226
rect 458138 496170 488678 496226
rect 488734 496170 488802 496226
rect 488858 496170 519398 496226
rect 519454 496170 519522 496226
rect 519578 496170 550118 496226
rect 550174 496170 550242 496226
rect 550298 496170 592914 496226
rect 592970 496170 593038 496226
rect 593094 496170 593162 496226
rect 593218 496170 593286 496226
rect 593342 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect -1916 496102 597980 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 27878 496102
rect 27934 496046 28002 496102
rect 28058 496046 58598 496102
rect 58654 496046 58722 496102
rect 58778 496046 89318 496102
rect 89374 496046 89442 496102
rect 89498 496046 120038 496102
rect 120094 496046 120162 496102
rect 120218 496046 150758 496102
rect 150814 496046 150882 496102
rect 150938 496046 181478 496102
rect 181534 496046 181602 496102
rect 181658 496046 212198 496102
rect 212254 496046 212322 496102
rect 212378 496046 242918 496102
rect 242974 496046 243042 496102
rect 243098 496046 273638 496102
rect 273694 496046 273762 496102
rect 273818 496046 304358 496102
rect 304414 496046 304482 496102
rect 304538 496046 335078 496102
rect 335134 496046 335202 496102
rect 335258 496046 365798 496102
rect 365854 496046 365922 496102
rect 365978 496046 396518 496102
rect 396574 496046 396642 496102
rect 396698 496046 427238 496102
rect 427294 496046 427362 496102
rect 427418 496046 457958 496102
rect 458014 496046 458082 496102
rect 458138 496046 488678 496102
rect 488734 496046 488802 496102
rect 488858 496046 519398 496102
rect 519454 496046 519522 496102
rect 519578 496046 550118 496102
rect 550174 496046 550242 496102
rect 550298 496046 592914 496102
rect 592970 496046 593038 496102
rect 593094 496046 593162 496102
rect 593218 496046 593286 496102
rect 593342 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect -1916 495978 597980 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 27878 495978
rect 27934 495922 28002 495978
rect 28058 495922 58598 495978
rect 58654 495922 58722 495978
rect 58778 495922 89318 495978
rect 89374 495922 89442 495978
rect 89498 495922 120038 495978
rect 120094 495922 120162 495978
rect 120218 495922 150758 495978
rect 150814 495922 150882 495978
rect 150938 495922 181478 495978
rect 181534 495922 181602 495978
rect 181658 495922 212198 495978
rect 212254 495922 212322 495978
rect 212378 495922 242918 495978
rect 242974 495922 243042 495978
rect 243098 495922 273638 495978
rect 273694 495922 273762 495978
rect 273818 495922 304358 495978
rect 304414 495922 304482 495978
rect 304538 495922 335078 495978
rect 335134 495922 335202 495978
rect 335258 495922 365798 495978
rect 365854 495922 365922 495978
rect 365978 495922 396518 495978
rect 396574 495922 396642 495978
rect 396698 495922 427238 495978
rect 427294 495922 427362 495978
rect 427418 495922 457958 495978
rect 458014 495922 458082 495978
rect 458138 495922 488678 495978
rect 488734 495922 488802 495978
rect 488858 495922 519398 495978
rect 519454 495922 519522 495978
rect 519578 495922 550118 495978
rect 550174 495922 550242 495978
rect 550298 495922 592914 495978
rect 592970 495922 593038 495978
rect 593094 495922 593162 495978
rect 593218 495922 593286 495978
rect 593342 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect -1916 495826 597980 495922
rect -1916 490350 597980 490446
rect -1916 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 5514 490350
rect 5570 490294 5638 490350
rect 5694 490294 5762 490350
rect 5818 490294 5886 490350
rect 5942 490294 12518 490350
rect 12574 490294 12642 490350
rect 12698 490294 43238 490350
rect 43294 490294 43362 490350
rect 43418 490294 73958 490350
rect 74014 490294 74082 490350
rect 74138 490294 104678 490350
rect 104734 490294 104802 490350
rect 104858 490294 135398 490350
rect 135454 490294 135522 490350
rect 135578 490294 166118 490350
rect 166174 490294 166242 490350
rect 166298 490294 196838 490350
rect 196894 490294 196962 490350
rect 197018 490294 227558 490350
rect 227614 490294 227682 490350
rect 227738 490294 258278 490350
rect 258334 490294 258402 490350
rect 258458 490294 288998 490350
rect 289054 490294 289122 490350
rect 289178 490294 319718 490350
rect 319774 490294 319842 490350
rect 319898 490294 350438 490350
rect 350494 490294 350562 490350
rect 350618 490294 381158 490350
rect 381214 490294 381282 490350
rect 381338 490294 411878 490350
rect 411934 490294 412002 490350
rect 412058 490294 442598 490350
rect 442654 490294 442722 490350
rect 442778 490294 473318 490350
rect 473374 490294 473442 490350
rect 473498 490294 504038 490350
rect 504094 490294 504162 490350
rect 504218 490294 534758 490350
rect 534814 490294 534882 490350
rect 534938 490294 565478 490350
rect 565534 490294 565602 490350
rect 565658 490294 589194 490350
rect 589250 490294 589318 490350
rect 589374 490294 589442 490350
rect 589498 490294 589566 490350
rect 589622 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597980 490350
rect -1916 490226 597980 490294
rect -1916 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 5514 490226
rect 5570 490170 5638 490226
rect 5694 490170 5762 490226
rect 5818 490170 5886 490226
rect 5942 490170 12518 490226
rect 12574 490170 12642 490226
rect 12698 490170 43238 490226
rect 43294 490170 43362 490226
rect 43418 490170 73958 490226
rect 74014 490170 74082 490226
rect 74138 490170 104678 490226
rect 104734 490170 104802 490226
rect 104858 490170 135398 490226
rect 135454 490170 135522 490226
rect 135578 490170 166118 490226
rect 166174 490170 166242 490226
rect 166298 490170 196838 490226
rect 196894 490170 196962 490226
rect 197018 490170 227558 490226
rect 227614 490170 227682 490226
rect 227738 490170 258278 490226
rect 258334 490170 258402 490226
rect 258458 490170 288998 490226
rect 289054 490170 289122 490226
rect 289178 490170 319718 490226
rect 319774 490170 319842 490226
rect 319898 490170 350438 490226
rect 350494 490170 350562 490226
rect 350618 490170 381158 490226
rect 381214 490170 381282 490226
rect 381338 490170 411878 490226
rect 411934 490170 412002 490226
rect 412058 490170 442598 490226
rect 442654 490170 442722 490226
rect 442778 490170 473318 490226
rect 473374 490170 473442 490226
rect 473498 490170 504038 490226
rect 504094 490170 504162 490226
rect 504218 490170 534758 490226
rect 534814 490170 534882 490226
rect 534938 490170 565478 490226
rect 565534 490170 565602 490226
rect 565658 490170 589194 490226
rect 589250 490170 589318 490226
rect 589374 490170 589442 490226
rect 589498 490170 589566 490226
rect 589622 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597980 490226
rect -1916 490102 597980 490170
rect -1916 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 5514 490102
rect 5570 490046 5638 490102
rect 5694 490046 5762 490102
rect 5818 490046 5886 490102
rect 5942 490046 12518 490102
rect 12574 490046 12642 490102
rect 12698 490046 43238 490102
rect 43294 490046 43362 490102
rect 43418 490046 73958 490102
rect 74014 490046 74082 490102
rect 74138 490046 104678 490102
rect 104734 490046 104802 490102
rect 104858 490046 135398 490102
rect 135454 490046 135522 490102
rect 135578 490046 166118 490102
rect 166174 490046 166242 490102
rect 166298 490046 196838 490102
rect 196894 490046 196962 490102
rect 197018 490046 227558 490102
rect 227614 490046 227682 490102
rect 227738 490046 258278 490102
rect 258334 490046 258402 490102
rect 258458 490046 288998 490102
rect 289054 490046 289122 490102
rect 289178 490046 319718 490102
rect 319774 490046 319842 490102
rect 319898 490046 350438 490102
rect 350494 490046 350562 490102
rect 350618 490046 381158 490102
rect 381214 490046 381282 490102
rect 381338 490046 411878 490102
rect 411934 490046 412002 490102
rect 412058 490046 442598 490102
rect 442654 490046 442722 490102
rect 442778 490046 473318 490102
rect 473374 490046 473442 490102
rect 473498 490046 504038 490102
rect 504094 490046 504162 490102
rect 504218 490046 534758 490102
rect 534814 490046 534882 490102
rect 534938 490046 565478 490102
rect 565534 490046 565602 490102
rect 565658 490046 589194 490102
rect 589250 490046 589318 490102
rect 589374 490046 589442 490102
rect 589498 490046 589566 490102
rect 589622 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597980 490102
rect -1916 489978 597980 490046
rect -1916 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 5514 489978
rect 5570 489922 5638 489978
rect 5694 489922 5762 489978
rect 5818 489922 5886 489978
rect 5942 489922 12518 489978
rect 12574 489922 12642 489978
rect 12698 489922 43238 489978
rect 43294 489922 43362 489978
rect 43418 489922 73958 489978
rect 74014 489922 74082 489978
rect 74138 489922 104678 489978
rect 104734 489922 104802 489978
rect 104858 489922 135398 489978
rect 135454 489922 135522 489978
rect 135578 489922 166118 489978
rect 166174 489922 166242 489978
rect 166298 489922 196838 489978
rect 196894 489922 196962 489978
rect 197018 489922 227558 489978
rect 227614 489922 227682 489978
rect 227738 489922 258278 489978
rect 258334 489922 258402 489978
rect 258458 489922 288998 489978
rect 289054 489922 289122 489978
rect 289178 489922 319718 489978
rect 319774 489922 319842 489978
rect 319898 489922 350438 489978
rect 350494 489922 350562 489978
rect 350618 489922 381158 489978
rect 381214 489922 381282 489978
rect 381338 489922 411878 489978
rect 411934 489922 412002 489978
rect 412058 489922 442598 489978
rect 442654 489922 442722 489978
rect 442778 489922 473318 489978
rect 473374 489922 473442 489978
rect 473498 489922 504038 489978
rect 504094 489922 504162 489978
rect 504218 489922 534758 489978
rect 534814 489922 534882 489978
rect 534938 489922 565478 489978
rect 565534 489922 565602 489978
rect 565658 489922 589194 489978
rect 589250 489922 589318 489978
rect 589374 489922 589442 489978
rect 589498 489922 589566 489978
rect 589622 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597980 489978
rect -1916 489826 597980 489922
rect -1916 478350 597980 478446
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 27878 478350
rect 27934 478294 28002 478350
rect 28058 478294 58598 478350
rect 58654 478294 58722 478350
rect 58778 478294 89318 478350
rect 89374 478294 89442 478350
rect 89498 478294 120038 478350
rect 120094 478294 120162 478350
rect 120218 478294 150758 478350
rect 150814 478294 150882 478350
rect 150938 478294 181478 478350
rect 181534 478294 181602 478350
rect 181658 478294 212198 478350
rect 212254 478294 212322 478350
rect 212378 478294 242918 478350
rect 242974 478294 243042 478350
rect 243098 478294 273638 478350
rect 273694 478294 273762 478350
rect 273818 478294 304358 478350
rect 304414 478294 304482 478350
rect 304538 478294 335078 478350
rect 335134 478294 335202 478350
rect 335258 478294 365798 478350
rect 365854 478294 365922 478350
rect 365978 478294 396518 478350
rect 396574 478294 396642 478350
rect 396698 478294 427238 478350
rect 427294 478294 427362 478350
rect 427418 478294 457958 478350
rect 458014 478294 458082 478350
rect 458138 478294 488678 478350
rect 488734 478294 488802 478350
rect 488858 478294 519398 478350
rect 519454 478294 519522 478350
rect 519578 478294 550118 478350
rect 550174 478294 550242 478350
rect 550298 478294 592914 478350
rect 592970 478294 593038 478350
rect 593094 478294 593162 478350
rect 593218 478294 593286 478350
rect 593342 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect -1916 478226 597980 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 27878 478226
rect 27934 478170 28002 478226
rect 28058 478170 58598 478226
rect 58654 478170 58722 478226
rect 58778 478170 89318 478226
rect 89374 478170 89442 478226
rect 89498 478170 120038 478226
rect 120094 478170 120162 478226
rect 120218 478170 150758 478226
rect 150814 478170 150882 478226
rect 150938 478170 181478 478226
rect 181534 478170 181602 478226
rect 181658 478170 212198 478226
rect 212254 478170 212322 478226
rect 212378 478170 242918 478226
rect 242974 478170 243042 478226
rect 243098 478170 273638 478226
rect 273694 478170 273762 478226
rect 273818 478170 304358 478226
rect 304414 478170 304482 478226
rect 304538 478170 335078 478226
rect 335134 478170 335202 478226
rect 335258 478170 365798 478226
rect 365854 478170 365922 478226
rect 365978 478170 396518 478226
rect 396574 478170 396642 478226
rect 396698 478170 427238 478226
rect 427294 478170 427362 478226
rect 427418 478170 457958 478226
rect 458014 478170 458082 478226
rect 458138 478170 488678 478226
rect 488734 478170 488802 478226
rect 488858 478170 519398 478226
rect 519454 478170 519522 478226
rect 519578 478170 550118 478226
rect 550174 478170 550242 478226
rect 550298 478170 592914 478226
rect 592970 478170 593038 478226
rect 593094 478170 593162 478226
rect 593218 478170 593286 478226
rect 593342 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect -1916 478102 597980 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 27878 478102
rect 27934 478046 28002 478102
rect 28058 478046 58598 478102
rect 58654 478046 58722 478102
rect 58778 478046 89318 478102
rect 89374 478046 89442 478102
rect 89498 478046 120038 478102
rect 120094 478046 120162 478102
rect 120218 478046 150758 478102
rect 150814 478046 150882 478102
rect 150938 478046 181478 478102
rect 181534 478046 181602 478102
rect 181658 478046 212198 478102
rect 212254 478046 212322 478102
rect 212378 478046 242918 478102
rect 242974 478046 243042 478102
rect 243098 478046 273638 478102
rect 273694 478046 273762 478102
rect 273818 478046 304358 478102
rect 304414 478046 304482 478102
rect 304538 478046 335078 478102
rect 335134 478046 335202 478102
rect 335258 478046 365798 478102
rect 365854 478046 365922 478102
rect 365978 478046 396518 478102
rect 396574 478046 396642 478102
rect 396698 478046 427238 478102
rect 427294 478046 427362 478102
rect 427418 478046 457958 478102
rect 458014 478046 458082 478102
rect 458138 478046 488678 478102
rect 488734 478046 488802 478102
rect 488858 478046 519398 478102
rect 519454 478046 519522 478102
rect 519578 478046 550118 478102
rect 550174 478046 550242 478102
rect 550298 478046 592914 478102
rect 592970 478046 593038 478102
rect 593094 478046 593162 478102
rect 593218 478046 593286 478102
rect 593342 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect -1916 477978 597980 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 27878 477978
rect 27934 477922 28002 477978
rect 28058 477922 58598 477978
rect 58654 477922 58722 477978
rect 58778 477922 89318 477978
rect 89374 477922 89442 477978
rect 89498 477922 120038 477978
rect 120094 477922 120162 477978
rect 120218 477922 150758 477978
rect 150814 477922 150882 477978
rect 150938 477922 181478 477978
rect 181534 477922 181602 477978
rect 181658 477922 212198 477978
rect 212254 477922 212322 477978
rect 212378 477922 242918 477978
rect 242974 477922 243042 477978
rect 243098 477922 273638 477978
rect 273694 477922 273762 477978
rect 273818 477922 304358 477978
rect 304414 477922 304482 477978
rect 304538 477922 335078 477978
rect 335134 477922 335202 477978
rect 335258 477922 365798 477978
rect 365854 477922 365922 477978
rect 365978 477922 396518 477978
rect 396574 477922 396642 477978
rect 396698 477922 427238 477978
rect 427294 477922 427362 477978
rect 427418 477922 457958 477978
rect 458014 477922 458082 477978
rect 458138 477922 488678 477978
rect 488734 477922 488802 477978
rect 488858 477922 519398 477978
rect 519454 477922 519522 477978
rect 519578 477922 550118 477978
rect 550174 477922 550242 477978
rect 550298 477922 592914 477978
rect 592970 477922 593038 477978
rect 593094 477922 593162 477978
rect 593218 477922 593286 477978
rect 593342 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect -1916 477826 597980 477922
rect -1916 472350 597980 472446
rect -1916 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 5514 472350
rect 5570 472294 5638 472350
rect 5694 472294 5762 472350
rect 5818 472294 5886 472350
rect 5942 472294 12518 472350
rect 12574 472294 12642 472350
rect 12698 472294 43238 472350
rect 43294 472294 43362 472350
rect 43418 472294 73958 472350
rect 74014 472294 74082 472350
rect 74138 472294 104678 472350
rect 104734 472294 104802 472350
rect 104858 472294 135398 472350
rect 135454 472294 135522 472350
rect 135578 472294 166118 472350
rect 166174 472294 166242 472350
rect 166298 472294 196838 472350
rect 196894 472294 196962 472350
rect 197018 472294 227558 472350
rect 227614 472294 227682 472350
rect 227738 472294 258278 472350
rect 258334 472294 258402 472350
rect 258458 472294 288998 472350
rect 289054 472294 289122 472350
rect 289178 472294 319718 472350
rect 319774 472294 319842 472350
rect 319898 472294 350438 472350
rect 350494 472294 350562 472350
rect 350618 472294 381158 472350
rect 381214 472294 381282 472350
rect 381338 472294 411878 472350
rect 411934 472294 412002 472350
rect 412058 472294 442598 472350
rect 442654 472294 442722 472350
rect 442778 472294 473318 472350
rect 473374 472294 473442 472350
rect 473498 472294 504038 472350
rect 504094 472294 504162 472350
rect 504218 472294 534758 472350
rect 534814 472294 534882 472350
rect 534938 472294 565478 472350
rect 565534 472294 565602 472350
rect 565658 472294 589194 472350
rect 589250 472294 589318 472350
rect 589374 472294 589442 472350
rect 589498 472294 589566 472350
rect 589622 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597980 472350
rect -1916 472226 597980 472294
rect -1916 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 5514 472226
rect 5570 472170 5638 472226
rect 5694 472170 5762 472226
rect 5818 472170 5886 472226
rect 5942 472170 12518 472226
rect 12574 472170 12642 472226
rect 12698 472170 43238 472226
rect 43294 472170 43362 472226
rect 43418 472170 73958 472226
rect 74014 472170 74082 472226
rect 74138 472170 104678 472226
rect 104734 472170 104802 472226
rect 104858 472170 135398 472226
rect 135454 472170 135522 472226
rect 135578 472170 166118 472226
rect 166174 472170 166242 472226
rect 166298 472170 196838 472226
rect 196894 472170 196962 472226
rect 197018 472170 227558 472226
rect 227614 472170 227682 472226
rect 227738 472170 258278 472226
rect 258334 472170 258402 472226
rect 258458 472170 288998 472226
rect 289054 472170 289122 472226
rect 289178 472170 319718 472226
rect 319774 472170 319842 472226
rect 319898 472170 350438 472226
rect 350494 472170 350562 472226
rect 350618 472170 381158 472226
rect 381214 472170 381282 472226
rect 381338 472170 411878 472226
rect 411934 472170 412002 472226
rect 412058 472170 442598 472226
rect 442654 472170 442722 472226
rect 442778 472170 473318 472226
rect 473374 472170 473442 472226
rect 473498 472170 504038 472226
rect 504094 472170 504162 472226
rect 504218 472170 534758 472226
rect 534814 472170 534882 472226
rect 534938 472170 565478 472226
rect 565534 472170 565602 472226
rect 565658 472170 589194 472226
rect 589250 472170 589318 472226
rect 589374 472170 589442 472226
rect 589498 472170 589566 472226
rect 589622 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597980 472226
rect -1916 472102 597980 472170
rect -1916 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 5514 472102
rect 5570 472046 5638 472102
rect 5694 472046 5762 472102
rect 5818 472046 5886 472102
rect 5942 472046 12518 472102
rect 12574 472046 12642 472102
rect 12698 472046 43238 472102
rect 43294 472046 43362 472102
rect 43418 472046 73958 472102
rect 74014 472046 74082 472102
rect 74138 472046 104678 472102
rect 104734 472046 104802 472102
rect 104858 472046 135398 472102
rect 135454 472046 135522 472102
rect 135578 472046 166118 472102
rect 166174 472046 166242 472102
rect 166298 472046 196838 472102
rect 196894 472046 196962 472102
rect 197018 472046 227558 472102
rect 227614 472046 227682 472102
rect 227738 472046 258278 472102
rect 258334 472046 258402 472102
rect 258458 472046 288998 472102
rect 289054 472046 289122 472102
rect 289178 472046 319718 472102
rect 319774 472046 319842 472102
rect 319898 472046 350438 472102
rect 350494 472046 350562 472102
rect 350618 472046 381158 472102
rect 381214 472046 381282 472102
rect 381338 472046 411878 472102
rect 411934 472046 412002 472102
rect 412058 472046 442598 472102
rect 442654 472046 442722 472102
rect 442778 472046 473318 472102
rect 473374 472046 473442 472102
rect 473498 472046 504038 472102
rect 504094 472046 504162 472102
rect 504218 472046 534758 472102
rect 534814 472046 534882 472102
rect 534938 472046 565478 472102
rect 565534 472046 565602 472102
rect 565658 472046 589194 472102
rect 589250 472046 589318 472102
rect 589374 472046 589442 472102
rect 589498 472046 589566 472102
rect 589622 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597980 472102
rect -1916 471978 597980 472046
rect -1916 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 5514 471978
rect 5570 471922 5638 471978
rect 5694 471922 5762 471978
rect 5818 471922 5886 471978
rect 5942 471922 12518 471978
rect 12574 471922 12642 471978
rect 12698 471922 43238 471978
rect 43294 471922 43362 471978
rect 43418 471922 73958 471978
rect 74014 471922 74082 471978
rect 74138 471922 104678 471978
rect 104734 471922 104802 471978
rect 104858 471922 135398 471978
rect 135454 471922 135522 471978
rect 135578 471922 166118 471978
rect 166174 471922 166242 471978
rect 166298 471922 196838 471978
rect 196894 471922 196962 471978
rect 197018 471922 227558 471978
rect 227614 471922 227682 471978
rect 227738 471922 258278 471978
rect 258334 471922 258402 471978
rect 258458 471922 288998 471978
rect 289054 471922 289122 471978
rect 289178 471922 319718 471978
rect 319774 471922 319842 471978
rect 319898 471922 350438 471978
rect 350494 471922 350562 471978
rect 350618 471922 381158 471978
rect 381214 471922 381282 471978
rect 381338 471922 411878 471978
rect 411934 471922 412002 471978
rect 412058 471922 442598 471978
rect 442654 471922 442722 471978
rect 442778 471922 473318 471978
rect 473374 471922 473442 471978
rect 473498 471922 504038 471978
rect 504094 471922 504162 471978
rect 504218 471922 534758 471978
rect 534814 471922 534882 471978
rect 534938 471922 565478 471978
rect 565534 471922 565602 471978
rect 565658 471922 589194 471978
rect 589250 471922 589318 471978
rect 589374 471922 589442 471978
rect 589498 471922 589566 471978
rect 589622 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597980 471978
rect -1916 471826 597980 471922
rect -1916 460350 597980 460446
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 27878 460350
rect 27934 460294 28002 460350
rect 28058 460294 58598 460350
rect 58654 460294 58722 460350
rect 58778 460294 89318 460350
rect 89374 460294 89442 460350
rect 89498 460294 120038 460350
rect 120094 460294 120162 460350
rect 120218 460294 150758 460350
rect 150814 460294 150882 460350
rect 150938 460294 181478 460350
rect 181534 460294 181602 460350
rect 181658 460294 212198 460350
rect 212254 460294 212322 460350
rect 212378 460294 242918 460350
rect 242974 460294 243042 460350
rect 243098 460294 273638 460350
rect 273694 460294 273762 460350
rect 273818 460294 304358 460350
rect 304414 460294 304482 460350
rect 304538 460294 335078 460350
rect 335134 460294 335202 460350
rect 335258 460294 365798 460350
rect 365854 460294 365922 460350
rect 365978 460294 396518 460350
rect 396574 460294 396642 460350
rect 396698 460294 427238 460350
rect 427294 460294 427362 460350
rect 427418 460294 457958 460350
rect 458014 460294 458082 460350
rect 458138 460294 488678 460350
rect 488734 460294 488802 460350
rect 488858 460294 519398 460350
rect 519454 460294 519522 460350
rect 519578 460294 550118 460350
rect 550174 460294 550242 460350
rect 550298 460294 592914 460350
rect 592970 460294 593038 460350
rect 593094 460294 593162 460350
rect 593218 460294 593286 460350
rect 593342 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect -1916 460226 597980 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 27878 460226
rect 27934 460170 28002 460226
rect 28058 460170 58598 460226
rect 58654 460170 58722 460226
rect 58778 460170 89318 460226
rect 89374 460170 89442 460226
rect 89498 460170 120038 460226
rect 120094 460170 120162 460226
rect 120218 460170 150758 460226
rect 150814 460170 150882 460226
rect 150938 460170 181478 460226
rect 181534 460170 181602 460226
rect 181658 460170 212198 460226
rect 212254 460170 212322 460226
rect 212378 460170 242918 460226
rect 242974 460170 243042 460226
rect 243098 460170 273638 460226
rect 273694 460170 273762 460226
rect 273818 460170 304358 460226
rect 304414 460170 304482 460226
rect 304538 460170 335078 460226
rect 335134 460170 335202 460226
rect 335258 460170 365798 460226
rect 365854 460170 365922 460226
rect 365978 460170 396518 460226
rect 396574 460170 396642 460226
rect 396698 460170 427238 460226
rect 427294 460170 427362 460226
rect 427418 460170 457958 460226
rect 458014 460170 458082 460226
rect 458138 460170 488678 460226
rect 488734 460170 488802 460226
rect 488858 460170 519398 460226
rect 519454 460170 519522 460226
rect 519578 460170 550118 460226
rect 550174 460170 550242 460226
rect 550298 460170 592914 460226
rect 592970 460170 593038 460226
rect 593094 460170 593162 460226
rect 593218 460170 593286 460226
rect 593342 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect -1916 460102 597980 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 27878 460102
rect 27934 460046 28002 460102
rect 28058 460046 58598 460102
rect 58654 460046 58722 460102
rect 58778 460046 89318 460102
rect 89374 460046 89442 460102
rect 89498 460046 120038 460102
rect 120094 460046 120162 460102
rect 120218 460046 150758 460102
rect 150814 460046 150882 460102
rect 150938 460046 181478 460102
rect 181534 460046 181602 460102
rect 181658 460046 212198 460102
rect 212254 460046 212322 460102
rect 212378 460046 242918 460102
rect 242974 460046 243042 460102
rect 243098 460046 273638 460102
rect 273694 460046 273762 460102
rect 273818 460046 304358 460102
rect 304414 460046 304482 460102
rect 304538 460046 335078 460102
rect 335134 460046 335202 460102
rect 335258 460046 365798 460102
rect 365854 460046 365922 460102
rect 365978 460046 396518 460102
rect 396574 460046 396642 460102
rect 396698 460046 427238 460102
rect 427294 460046 427362 460102
rect 427418 460046 457958 460102
rect 458014 460046 458082 460102
rect 458138 460046 488678 460102
rect 488734 460046 488802 460102
rect 488858 460046 519398 460102
rect 519454 460046 519522 460102
rect 519578 460046 550118 460102
rect 550174 460046 550242 460102
rect 550298 460046 592914 460102
rect 592970 460046 593038 460102
rect 593094 460046 593162 460102
rect 593218 460046 593286 460102
rect 593342 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect -1916 459978 597980 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 27878 459978
rect 27934 459922 28002 459978
rect 28058 459922 58598 459978
rect 58654 459922 58722 459978
rect 58778 459922 89318 459978
rect 89374 459922 89442 459978
rect 89498 459922 120038 459978
rect 120094 459922 120162 459978
rect 120218 459922 150758 459978
rect 150814 459922 150882 459978
rect 150938 459922 181478 459978
rect 181534 459922 181602 459978
rect 181658 459922 212198 459978
rect 212254 459922 212322 459978
rect 212378 459922 242918 459978
rect 242974 459922 243042 459978
rect 243098 459922 273638 459978
rect 273694 459922 273762 459978
rect 273818 459922 304358 459978
rect 304414 459922 304482 459978
rect 304538 459922 335078 459978
rect 335134 459922 335202 459978
rect 335258 459922 365798 459978
rect 365854 459922 365922 459978
rect 365978 459922 396518 459978
rect 396574 459922 396642 459978
rect 396698 459922 427238 459978
rect 427294 459922 427362 459978
rect 427418 459922 457958 459978
rect 458014 459922 458082 459978
rect 458138 459922 488678 459978
rect 488734 459922 488802 459978
rect 488858 459922 519398 459978
rect 519454 459922 519522 459978
rect 519578 459922 550118 459978
rect 550174 459922 550242 459978
rect 550298 459922 592914 459978
rect 592970 459922 593038 459978
rect 593094 459922 593162 459978
rect 593218 459922 593286 459978
rect 593342 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect -1916 459826 597980 459922
rect -1916 454350 597980 454446
rect -1916 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 5514 454350
rect 5570 454294 5638 454350
rect 5694 454294 5762 454350
rect 5818 454294 5886 454350
rect 5942 454294 12518 454350
rect 12574 454294 12642 454350
rect 12698 454294 43238 454350
rect 43294 454294 43362 454350
rect 43418 454294 73958 454350
rect 74014 454294 74082 454350
rect 74138 454294 104678 454350
rect 104734 454294 104802 454350
rect 104858 454294 135398 454350
rect 135454 454294 135522 454350
rect 135578 454294 166118 454350
rect 166174 454294 166242 454350
rect 166298 454294 196838 454350
rect 196894 454294 196962 454350
rect 197018 454294 227558 454350
rect 227614 454294 227682 454350
rect 227738 454294 258278 454350
rect 258334 454294 258402 454350
rect 258458 454294 288998 454350
rect 289054 454294 289122 454350
rect 289178 454294 319718 454350
rect 319774 454294 319842 454350
rect 319898 454294 350438 454350
rect 350494 454294 350562 454350
rect 350618 454294 381158 454350
rect 381214 454294 381282 454350
rect 381338 454294 411878 454350
rect 411934 454294 412002 454350
rect 412058 454294 442598 454350
rect 442654 454294 442722 454350
rect 442778 454294 473318 454350
rect 473374 454294 473442 454350
rect 473498 454294 504038 454350
rect 504094 454294 504162 454350
rect 504218 454294 534758 454350
rect 534814 454294 534882 454350
rect 534938 454294 565478 454350
rect 565534 454294 565602 454350
rect 565658 454294 589194 454350
rect 589250 454294 589318 454350
rect 589374 454294 589442 454350
rect 589498 454294 589566 454350
rect 589622 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597980 454350
rect -1916 454226 597980 454294
rect -1916 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 5514 454226
rect 5570 454170 5638 454226
rect 5694 454170 5762 454226
rect 5818 454170 5886 454226
rect 5942 454170 12518 454226
rect 12574 454170 12642 454226
rect 12698 454170 43238 454226
rect 43294 454170 43362 454226
rect 43418 454170 73958 454226
rect 74014 454170 74082 454226
rect 74138 454170 104678 454226
rect 104734 454170 104802 454226
rect 104858 454170 135398 454226
rect 135454 454170 135522 454226
rect 135578 454170 166118 454226
rect 166174 454170 166242 454226
rect 166298 454170 196838 454226
rect 196894 454170 196962 454226
rect 197018 454170 227558 454226
rect 227614 454170 227682 454226
rect 227738 454170 258278 454226
rect 258334 454170 258402 454226
rect 258458 454170 288998 454226
rect 289054 454170 289122 454226
rect 289178 454170 319718 454226
rect 319774 454170 319842 454226
rect 319898 454170 350438 454226
rect 350494 454170 350562 454226
rect 350618 454170 381158 454226
rect 381214 454170 381282 454226
rect 381338 454170 411878 454226
rect 411934 454170 412002 454226
rect 412058 454170 442598 454226
rect 442654 454170 442722 454226
rect 442778 454170 473318 454226
rect 473374 454170 473442 454226
rect 473498 454170 504038 454226
rect 504094 454170 504162 454226
rect 504218 454170 534758 454226
rect 534814 454170 534882 454226
rect 534938 454170 565478 454226
rect 565534 454170 565602 454226
rect 565658 454170 589194 454226
rect 589250 454170 589318 454226
rect 589374 454170 589442 454226
rect 589498 454170 589566 454226
rect 589622 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597980 454226
rect -1916 454102 597980 454170
rect -1916 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 5514 454102
rect 5570 454046 5638 454102
rect 5694 454046 5762 454102
rect 5818 454046 5886 454102
rect 5942 454046 12518 454102
rect 12574 454046 12642 454102
rect 12698 454046 43238 454102
rect 43294 454046 43362 454102
rect 43418 454046 73958 454102
rect 74014 454046 74082 454102
rect 74138 454046 104678 454102
rect 104734 454046 104802 454102
rect 104858 454046 135398 454102
rect 135454 454046 135522 454102
rect 135578 454046 166118 454102
rect 166174 454046 166242 454102
rect 166298 454046 196838 454102
rect 196894 454046 196962 454102
rect 197018 454046 227558 454102
rect 227614 454046 227682 454102
rect 227738 454046 258278 454102
rect 258334 454046 258402 454102
rect 258458 454046 288998 454102
rect 289054 454046 289122 454102
rect 289178 454046 319718 454102
rect 319774 454046 319842 454102
rect 319898 454046 350438 454102
rect 350494 454046 350562 454102
rect 350618 454046 381158 454102
rect 381214 454046 381282 454102
rect 381338 454046 411878 454102
rect 411934 454046 412002 454102
rect 412058 454046 442598 454102
rect 442654 454046 442722 454102
rect 442778 454046 473318 454102
rect 473374 454046 473442 454102
rect 473498 454046 504038 454102
rect 504094 454046 504162 454102
rect 504218 454046 534758 454102
rect 534814 454046 534882 454102
rect 534938 454046 565478 454102
rect 565534 454046 565602 454102
rect 565658 454046 589194 454102
rect 589250 454046 589318 454102
rect 589374 454046 589442 454102
rect 589498 454046 589566 454102
rect 589622 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597980 454102
rect -1916 453978 597980 454046
rect -1916 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 5514 453978
rect 5570 453922 5638 453978
rect 5694 453922 5762 453978
rect 5818 453922 5886 453978
rect 5942 453922 12518 453978
rect 12574 453922 12642 453978
rect 12698 453922 43238 453978
rect 43294 453922 43362 453978
rect 43418 453922 73958 453978
rect 74014 453922 74082 453978
rect 74138 453922 104678 453978
rect 104734 453922 104802 453978
rect 104858 453922 135398 453978
rect 135454 453922 135522 453978
rect 135578 453922 166118 453978
rect 166174 453922 166242 453978
rect 166298 453922 196838 453978
rect 196894 453922 196962 453978
rect 197018 453922 227558 453978
rect 227614 453922 227682 453978
rect 227738 453922 258278 453978
rect 258334 453922 258402 453978
rect 258458 453922 288998 453978
rect 289054 453922 289122 453978
rect 289178 453922 319718 453978
rect 319774 453922 319842 453978
rect 319898 453922 350438 453978
rect 350494 453922 350562 453978
rect 350618 453922 381158 453978
rect 381214 453922 381282 453978
rect 381338 453922 411878 453978
rect 411934 453922 412002 453978
rect 412058 453922 442598 453978
rect 442654 453922 442722 453978
rect 442778 453922 473318 453978
rect 473374 453922 473442 453978
rect 473498 453922 504038 453978
rect 504094 453922 504162 453978
rect 504218 453922 534758 453978
rect 534814 453922 534882 453978
rect 534938 453922 565478 453978
rect 565534 453922 565602 453978
rect 565658 453922 589194 453978
rect 589250 453922 589318 453978
rect 589374 453922 589442 453978
rect 589498 453922 589566 453978
rect 589622 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597980 453978
rect -1916 453826 597980 453922
rect -1916 442350 597980 442446
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 27878 442350
rect 27934 442294 28002 442350
rect 28058 442294 58598 442350
rect 58654 442294 58722 442350
rect 58778 442294 89318 442350
rect 89374 442294 89442 442350
rect 89498 442294 120038 442350
rect 120094 442294 120162 442350
rect 120218 442294 150758 442350
rect 150814 442294 150882 442350
rect 150938 442294 181478 442350
rect 181534 442294 181602 442350
rect 181658 442294 212198 442350
rect 212254 442294 212322 442350
rect 212378 442294 242918 442350
rect 242974 442294 243042 442350
rect 243098 442294 273638 442350
rect 273694 442294 273762 442350
rect 273818 442294 304358 442350
rect 304414 442294 304482 442350
rect 304538 442294 335078 442350
rect 335134 442294 335202 442350
rect 335258 442294 365798 442350
rect 365854 442294 365922 442350
rect 365978 442294 396518 442350
rect 396574 442294 396642 442350
rect 396698 442294 427238 442350
rect 427294 442294 427362 442350
rect 427418 442294 457958 442350
rect 458014 442294 458082 442350
rect 458138 442294 488678 442350
rect 488734 442294 488802 442350
rect 488858 442294 519398 442350
rect 519454 442294 519522 442350
rect 519578 442294 550118 442350
rect 550174 442294 550242 442350
rect 550298 442294 592914 442350
rect 592970 442294 593038 442350
rect 593094 442294 593162 442350
rect 593218 442294 593286 442350
rect 593342 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect -1916 442226 597980 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 27878 442226
rect 27934 442170 28002 442226
rect 28058 442170 58598 442226
rect 58654 442170 58722 442226
rect 58778 442170 89318 442226
rect 89374 442170 89442 442226
rect 89498 442170 120038 442226
rect 120094 442170 120162 442226
rect 120218 442170 150758 442226
rect 150814 442170 150882 442226
rect 150938 442170 181478 442226
rect 181534 442170 181602 442226
rect 181658 442170 212198 442226
rect 212254 442170 212322 442226
rect 212378 442170 242918 442226
rect 242974 442170 243042 442226
rect 243098 442170 273638 442226
rect 273694 442170 273762 442226
rect 273818 442170 304358 442226
rect 304414 442170 304482 442226
rect 304538 442170 335078 442226
rect 335134 442170 335202 442226
rect 335258 442170 365798 442226
rect 365854 442170 365922 442226
rect 365978 442170 396518 442226
rect 396574 442170 396642 442226
rect 396698 442170 427238 442226
rect 427294 442170 427362 442226
rect 427418 442170 457958 442226
rect 458014 442170 458082 442226
rect 458138 442170 488678 442226
rect 488734 442170 488802 442226
rect 488858 442170 519398 442226
rect 519454 442170 519522 442226
rect 519578 442170 550118 442226
rect 550174 442170 550242 442226
rect 550298 442170 592914 442226
rect 592970 442170 593038 442226
rect 593094 442170 593162 442226
rect 593218 442170 593286 442226
rect 593342 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect -1916 442102 597980 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 27878 442102
rect 27934 442046 28002 442102
rect 28058 442046 58598 442102
rect 58654 442046 58722 442102
rect 58778 442046 89318 442102
rect 89374 442046 89442 442102
rect 89498 442046 120038 442102
rect 120094 442046 120162 442102
rect 120218 442046 150758 442102
rect 150814 442046 150882 442102
rect 150938 442046 181478 442102
rect 181534 442046 181602 442102
rect 181658 442046 212198 442102
rect 212254 442046 212322 442102
rect 212378 442046 242918 442102
rect 242974 442046 243042 442102
rect 243098 442046 273638 442102
rect 273694 442046 273762 442102
rect 273818 442046 304358 442102
rect 304414 442046 304482 442102
rect 304538 442046 335078 442102
rect 335134 442046 335202 442102
rect 335258 442046 365798 442102
rect 365854 442046 365922 442102
rect 365978 442046 396518 442102
rect 396574 442046 396642 442102
rect 396698 442046 427238 442102
rect 427294 442046 427362 442102
rect 427418 442046 457958 442102
rect 458014 442046 458082 442102
rect 458138 442046 488678 442102
rect 488734 442046 488802 442102
rect 488858 442046 519398 442102
rect 519454 442046 519522 442102
rect 519578 442046 550118 442102
rect 550174 442046 550242 442102
rect 550298 442046 592914 442102
rect 592970 442046 593038 442102
rect 593094 442046 593162 442102
rect 593218 442046 593286 442102
rect 593342 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect -1916 441978 597980 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 27878 441978
rect 27934 441922 28002 441978
rect 28058 441922 58598 441978
rect 58654 441922 58722 441978
rect 58778 441922 89318 441978
rect 89374 441922 89442 441978
rect 89498 441922 120038 441978
rect 120094 441922 120162 441978
rect 120218 441922 150758 441978
rect 150814 441922 150882 441978
rect 150938 441922 181478 441978
rect 181534 441922 181602 441978
rect 181658 441922 212198 441978
rect 212254 441922 212322 441978
rect 212378 441922 242918 441978
rect 242974 441922 243042 441978
rect 243098 441922 273638 441978
rect 273694 441922 273762 441978
rect 273818 441922 304358 441978
rect 304414 441922 304482 441978
rect 304538 441922 335078 441978
rect 335134 441922 335202 441978
rect 335258 441922 365798 441978
rect 365854 441922 365922 441978
rect 365978 441922 396518 441978
rect 396574 441922 396642 441978
rect 396698 441922 427238 441978
rect 427294 441922 427362 441978
rect 427418 441922 457958 441978
rect 458014 441922 458082 441978
rect 458138 441922 488678 441978
rect 488734 441922 488802 441978
rect 488858 441922 519398 441978
rect 519454 441922 519522 441978
rect 519578 441922 550118 441978
rect 550174 441922 550242 441978
rect 550298 441922 592914 441978
rect 592970 441922 593038 441978
rect 593094 441922 593162 441978
rect 593218 441922 593286 441978
rect 593342 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect -1916 441826 597980 441922
rect -1916 436350 597980 436446
rect -1916 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 5514 436350
rect 5570 436294 5638 436350
rect 5694 436294 5762 436350
rect 5818 436294 5886 436350
rect 5942 436294 12518 436350
rect 12574 436294 12642 436350
rect 12698 436294 43238 436350
rect 43294 436294 43362 436350
rect 43418 436294 73958 436350
rect 74014 436294 74082 436350
rect 74138 436294 104678 436350
rect 104734 436294 104802 436350
rect 104858 436294 135398 436350
rect 135454 436294 135522 436350
rect 135578 436294 166118 436350
rect 166174 436294 166242 436350
rect 166298 436294 196838 436350
rect 196894 436294 196962 436350
rect 197018 436294 227558 436350
rect 227614 436294 227682 436350
rect 227738 436294 258278 436350
rect 258334 436294 258402 436350
rect 258458 436294 288998 436350
rect 289054 436294 289122 436350
rect 289178 436294 319718 436350
rect 319774 436294 319842 436350
rect 319898 436294 350438 436350
rect 350494 436294 350562 436350
rect 350618 436294 381158 436350
rect 381214 436294 381282 436350
rect 381338 436294 411878 436350
rect 411934 436294 412002 436350
rect 412058 436294 442598 436350
rect 442654 436294 442722 436350
rect 442778 436294 473318 436350
rect 473374 436294 473442 436350
rect 473498 436294 504038 436350
rect 504094 436294 504162 436350
rect 504218 436294 534758 436350
rect 534814 436294 534882 436350
rect 534938 436294 565478 436350
rect 565534 436294 565602 436350
rect 565658 436294 589194 436350
rect 589250 436294 589318 436350
rect 589374 436294 589442 436350
rect 589498 436294 589566 436350
rect 589622 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597980 436350
rect -1916 436226 597980 436294
rect -1916 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 5514 436226
rect 5570 436170 5638 436226
rect 5694 436170 5762 436226
rect 5818 436170 5886 436226
rect 5942 436170 12518 436226
rect 12574 436170 12642 436226
rect 12698 436170 43238 436226
rect 43294 436170 43362 436226
rect 43418 436170 73958 436226
rect 74014 436170 74082 436226
rect 74138 436170 104678 436226
rect 104734 436170 104802 436226
rect 104858 436170 135398 436226
rect 135454 436170 135522 436226
rect 135578 436170 166118 436226
rect 166174 436170 166242 436226
rect 166298 436170 196838 436226
rect 196894 436170 196962 436226
rect 197018 436170 227558 436226
rect 227614 436170 227682 436226
rect 227738 436170 258278 436226
rect 258334 436170 258402 436226
rect 258458 436170 288998 436226
rect 289054 436170 289122 436226
rect 289178 436170 319718 436226
rect 319774 436170 319842 436226
rect 319898 436170 350438 436226
rect 350494 436170 350562 436226
rect 350618 436170 381158 436226
rect 381214 436170 381282 436226
rect 381338 436170 411878 436226
rect 411934 436170 412002 436226
rect 412058 436170 442598 436226
rect 442654 436170 442722 436226
rect 442778 436170 473318 436226
rect 473374 436170 473442 436226
rect 473498 436170 504038 436226
rect 504094 436170 504162 436226
rect 504218 436170 534758 436226
rect 534814 436170 534882 436226
rect 534938 436170 565478 436226
rect 565534 436170 565602 436226
rect 565658 436170 589194 436226
rect 589250 436170 589318 436226
rect 589374 436170 589442 436226
rect 589498 436170 589566 436226
rect 589622 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597980 436226
rect -1916 436102 597980 436170
rect -1916 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 5514 436102
rect 5570 436046 5638 436102
rect 5694 436046 5762 436102
rect 5818 436046 5886 436102
rect 5942 436046 12518 436102
rect 12574 436046 12642 436102
rect 12698 436046 43238 436102
rect 43294 436046 43362 436102
rect 43418 436046 73958 436102
rect 74014 436046 74082 436102
rect 74138 436046 104678 436102
rect 104734 436046 104802 436102
rect 104858 436046 135398 436102
rect 135454 436046 135522 436102
rect 135578 436046 166118 436102
rect 166174 436046 166242 436102
rect 166298 436046 196838 436102
rect 196894 436046 196962 436102
rect 197018 436046 227558 436102
rect 227614 436046 227682 436102
rect 227738 436046 258278 436102
rect 258334 436046 258402 436102
rect 258458 436046 288998 436102
rect 289054 436046 289122 436102
rect 289178 436046 319718 436102
rect 319774 436046 319842 436102
rect 319898 436046 350438 436102
rect 350494 436046 350562 436102
rect 350618 436046 381158 436102
rect 381214 436046 381282 436102
rect 381338 436046 411878 436102
rect 411934 436046 412002 436102
rect 412058 436046 442598 436102
rect 442654 436046 442722 436102
rect 442778 436046 473318 436102
rect 473374 436046 473442 436102
rect 473498 436046 504038 436102
rect 504094 436046 504162 436102
rect 504218 436046 534758 436102
rect 534814 436046 534882 436102
rect 534938 436046 565478 436102
rect 565534 436046 565602 436102
rect 565658 436046 589194 436102
rect 589250 436046 589318 436102
rect 589374 436046 589442 436102
rect 589498 436046 589566 436102
rect 589622 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597980 436102
rect -1916 435978 597980 436046
rect -1916 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 5514 435978
rect 5570 435922 5638 435978
rect 5694 435922 5762 435978
rect 5818 435922 5886 435978
rect 5942 435922 12518 435978
rect 12574 435922 12642 435978
rect 12698 435922 43238 435978
rect 43294 435922 43362 435978
rect 43418 435922 73958 435978
rect 74014 435922 74082 435978
rect 74138 435922 104678 435978
rect 104734 435922 104802 435978
rect 104858 435922 135398 435978
rect 135454 435922 135522 435978
rect 135578 435922 166118 435978
rect 166174 435922 166242 435978
rect 166298 435922 196838 435978
rect 196894 435922 196962 435978
rect 197018 435922 227558 435978
rect 227614 435922 227682 435978
rect 227738 435922 258278 435978
rect 258334 435922 258402 435978
rect 258458 435922 288998 435978
rect 289054 435922 289122 435978
rect 289178 435922 319718 435978
rect 319774 435922 319842 435978
rect 319898 435922 350438 435978
rect 350494 435922 350562 435978
rect 350618 435922 381158 435978
rect 381214 435922 381282 435978
rect 381338 435922 411878 435978
rect 411934 435922 412002 435978
rect 412058 435922 442598 435978
rect 442654 435922 442722 435978
rect 442778 435922 473318 435978
rect 473374 435922 473442 435978
rect 473498 435922 504038 435978
rect 504094 435922 504162 435978
rect 504218 435922 534758 435978
rect 534814 435922 534882 435978
rect 534938 435922 565478 435978
rect 565534 435922 565602 435978
rect 565658 435922 589194 435978
rect 589250 435922 589318 435978
rect 589374 435922 589442 435978
rect 589498 435922 589566 435978
rect 589622 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597980 435978
rect -1916 435826 597980 435922
rect -1916 424350 597980 424446
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 27878 424350
rect 27934 424294 28002 424350
rect 28058 424294 58598 424350
rect 58654 424294 58722 424350
rect 58778 424294 89318 424350
rect 89374 424294 89442 424350
rect 89498 424294 120038 424350
rect 120094 424294 120162 424350
rect 120218 424294 150758 424350
rect 150814 424294 150882 424350
rect 150938 424294 181478 424350
rect 181534 424294 181602 424350
rect 181658 424294 212198 424350
rect 212254 424294 212322 424350
rect 212378 424294 242918 424350
rect 242974 424294 243042 424350
rect 243098 424294 273638 424350
rect 273694 424294 273762 424350
rect 273818 424294 304358 424350
rect 304414 424294 304482 424350
rect 304538 424294 335078 424350
rect 335134 424294 335202 424350
rect 335258 424294 365798 424350
rect 365854 424294 365922 424350
rect 365978 424294 396518 424350
rect 396574 424294 396642 424350
rect 396698 424294 427238 424350
rect 427294 424294 427362 424350
rect 427418 424294 457958 424350
rect 458014 424294 458082 424350
rect 458138 424294 488678 424350
rect 488734 424294 488802 424350
rect 488858 424294 519398 424350
rect 519454 424294 519522 424350
rect 519578 424294 550118 424350
rect 550174 424294 550242 424350
rect 550298 424294 592914 424350
rect 592970 424294 593038 424350
rect 593094 424294 593162 424350
rect 593218 424294 593286 424350
rect 593342 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect -1916 424226 597980 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 27878 424226
rect 27934 424170 28002 424226
rect 28058 424170 58598 424226
rect 58654 424170 58722 424226
rect 58778 424170 89318 424226
rect 89374 424170 89442 424226
rect 89498 424170 120038 424226
rect 120094 424170 120162 424226
rect 120218 424170 150758 424226
rect 150814 424170 150882 424226
rect 150938 424170 181478 424226
rect 181534 424170 181602 424226
rect 181658 424170 212198 424226
rect 212254 424170 212322 424226
rect 212378 424170 242918 424226
rect 242974 424170 243042 424226
rect 243098 424170 273638 424226
rect 273694 424170 273762 424226
rect 273818 424170 304358 424226
rect 304414 424170 304482 424226
rect 304538 424170 335078 424226
rect 335134 424170 335202 424226
rect 335258 424170 365798 424226
rect 365854 424170 365922 424226
rect 365978 424170 396518 424226
rect 396574 424170 396642 424226
rect 396698 424170 427238 424226
rect 427294 424170 427362 424226
rect 427418 424170 457958 424226
rect 458014 424170 458082 424226
rect 458138 424170 488678 424226
rect 488734 424170 488802 424226
rect 488858 424170 519398 424226
rect 519454 424170 519522 424226
rect 519578 424170 550118 424226
rect 550174 424170 550242 424226
rect 550298 424170 592914 424226
rect 592970 424170 593038 424226
rect 593094 424170 593162 424226
rect 593218 424170 593286 424226
rect 593342 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect -1916 424102 597980 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 27878 424102
rect 27934 424046 28002 424102
rect 28058 424046 58598 424102
rect 58654 424046 58722 424102
rect 58778 424046 89318 424102
rect 89374 424046 89442 424102
rect 89498 424046 120038 424102
rect 120094 424046 120162 424102
rect 120218 424046 150758 424102
rect 150814 424046 150882 424102
rect 150938 424046 181478 424102
rect 181534 424046 181602 424102
rect 181658 424046 212198 424102
rect 212254 424046 212322 424102
rect 212378 424046 242918 424102
rect 242974 424046 243042 424102
rect 243098 424046 273638 424102
rect 273694 424046 273762 424102
rect 273818 424046 304358 424102
rect 304414 424046 304482 424102
rect 304538 424046 335078 424102
rect 335134 424046 335202 424102
rect 335258 424046 365798 424102
rect 365854 424046 365922 424102
rect 365978 424046 396518 424102
rect 396574 424046 396642 424102
rect 396698 424046 427238 424102
rect 427294 424046 427362 424102
rect 427418 424046 457958 424102
rect 458014 424046 458082 424102
rect 458138 424046 488678 424102
rect 488734 424046 488802 424102
rect 488858 424046 519398 424102
rect 519454 424046 519522 424102
rect 519578 424046 550118 424102
rect 550174 424046 550242 424102
rect 550298 424046 592914 424102
rect 592970 424046 593038 424102
rect 593094 424046 593162 424102
rect 593218 424046 593286 424102
rect 593342 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect -1916 423978 597980 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 27878 423978
rect 27934 423922 28002 423978
rect 28058 423922 58598 423978
rect 58654 423922 58722 423978
rect 58778 423922 89318 423978
rect 89374 423922 89442 423978
rect 89498 423922 120038 423978
rect 120094 423922 120162 423978
rect 120218 423922 150758 423978
rect 150814 423922 150882 423978
rect 150938 423922 181478 423978
rect 181534 423922 181602 423978
rect 181658 423922 212198 423978
rect 212254 423922 212322 423978
rect 212378 423922 242918 423978
rect 242974 423922 243042 423978
rect 243098 423922 273638 423978
rect 273694 423922 273762 423978
rect 273818 423922 304358 423978
rect 304414 423922 304482 423978
rect 304538 423922 335078 423978
rect 335134 423922 335202 423978
rect 335258 423922 365798 423978
rect 365854 423922 365922 423978
rect 365978 423922 396518 423978
rect 396574 423922 396642 423978
rect 396698 423922 427238 423978
rect 427294 423922 427362 423978
rect 427418 423922 457958 423978
rect 458014 423922 458082 423978
rect 458138 423922 488678 423978
rect 488734 423922 488802 423978
rect 488858 423922 519398 423978
rect 519454 423922 519522 423978
rect 519578 423922 550118 423978
rect 550174 423922 550242 423978
rect 550298 423922 592914 423978
rect 592970 423922 593038 423978
rect 593094 423922 593162 423978
rect 593218 423922 593286 423978
rect 593342 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect -1916 423826 597980 423922
rect -1916 418350 597980 418446
rect -1916 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 5514 418350
rect 5570 418294 5638 418350
rect 5694 418294 5762 418350
rect 5818 418294 5886 418350
rect 5942 418294 12518 418350
rect 12574 418294 12642 418350
rect 12698 418294 43238 418350
rect 43294 418294 43362 418350
rect 43418 418294 73958 418350
rect 74014 418294 74082 418350
rect 74138 418294 104678 418350
rect 104734 418294 104802 418350
rect 104858 418294 135398 418350
rect 135454 418294 135522 418350
rect 135578 418294 166118 418350
rect 166174 418294 166242 418350
rect 166298 418294 196838 418350
rect 196894 418294 196962 418350
rect 197018 418294 227558 418350
rect 227614 418294 227682 418350
rect 227738 418294 258278 418350
rect 258334 418294 258402 418350
rect 258458 418294 288998 418350
rect 289054 418294 289122 418350
rect 289178 418294 319718 418350
rect 319774 418294 319842 418350
rect 319898 418294 350438 418350
rect 350494 418294 350562 418350
rect 350618 418294 381158 418350
rect 381214 418294 381282 418350
rect 381338 418294 411878 418350
rect 411934 418294 412002 418350
rect 412058 418294 442598 418350
rect 442654 418294 442722 418350
rect 442778 418294 473318 418350
rect 473374 418294 473442 418350
rect 473498 418294 504038 418350
rect 504094 418294 504162 418350
rect 504218 418294 534758 418350
rect 534814 418294 534882 418350
rect 534938 418294 565478 418350
rect 565534 418294 565602 418350
rect 565658 418294 589194 418350
rect 589250 418294 589318 418350
rect 589374 418294 589442 418350
rect 589498 418294 589566 418350
rect 589622 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597980 418350
rect -1916 418226 597980 418294
rect -1916 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 5514 418226
rect 5570 418170 5638 418226
rect 5694 418170 5762 418226
rect 5818 418170 5886 418226
rect 5942 418170 12518 418226
rect 12574 418170 12642 418226
rect 12698 418170 43238 418226
rect 43294 418170 43362 418226
rect 43418 418170 73958 418226
rect 74014 418170 74082 418226
rect 74138 418170 104678 418226
rect 104734 418170 104802 418226
rect 104858 418170 135398 418226
rect 135454 418170 135522 418226
rect 135578 418170 166118 418226
rect 166174 418170 166242 418226
rect 166298 418170 196838 418226
rect 196894 418170 196962 418226
rect 197018 418170 227558 418226
rect 227614 418170 227682 418226
rect 227738 418170 258278 418226
rect 258334 418170 258402 418226
rect 258458 418170 288998 418226
rect 289054 418170 289122 418226
rect 289178 418170 319718 418226
rect 319774 418170 319842 418226
rect 319898 418170 350438 418226
rect 350494 418170 350562 418226
rect 350618 418170 381158 418226
rect 381214 418170 381282 418226
rect 381338 418170 411878 418226
rect 411934 418170 412002 418226
rect 412058 418170 442598 418226
rect 442654 418170 442722 418226
rect 442778 418170 473318 418226
rect 473374 418170 473442 418226
rect 473498 418170 504038 418226
rect 504094 418170 504162 418226
rect 504218 418170 534758 418226
rect 534814 418170 534882 418226
rect 534938 418170 565478 418226
rect 565534 418170 565602 418226
rect 565658 418170 589194 418226
rect 589250 418170 589318 418226
rect 589374 418170 589442 418226
rect 589498 418170 589566 418226
rect 589622 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597980 418226
rect -1916 418102 597980 418170
rect -1916 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 5514 418102
rect 5570 418046 5638 418102
rect 5694 418046 5762 418102
rect 5818 418046 5886 418102
rect 5942 418046 12518 418102
rect 12574 418046 12642 418102
rect 12698 418046 43238 418102
rect 43294 418046 43362 418102
rect 43418 418046 73958 418102
rect 74014 418046 74082 418102
rect 74138 418046 104678 418102
rect 104734 418046 104802 418102
rect 104858 418046 135398 418102
rect 135454 418046 135522 418102
rect 135578 418046 166118 418102
rect 166174 418046 166242 418102
rect 166298 418046 196838 418102
rect 196894 418046 196962 418102
rect 197018 418046 227558 418102
rect 227614 418046 227682 418102
rect 227738 418046 258278 418102
rect 258334 418046 258402 418102
rect 258458 418046 288998 418102
rect 289054 418046 289122 418102
rect 289178 418046 319718 418102
rect 319774 418046 319842 418102
rect 319898 418046 350438 418102
rect 350494 418046 350562 418102
rect 350618 418046 381158 418102
rect 381214 418046 381282 418102
rect 381338 418046 411878 418102
rect 411934 418046 412002 418102
rect 412058 418046 442598 418102
rect 442654 418046 442722 418102
rect 442778 418046 473318 418102
rect 473374 418046 473442 418102
rect 473498 418046 504038 418102
rect 504094 418046 504162 418102
rect 504218 418046 534758 418102
rect 534814 418046 534882 418102
rect 534938 418046 565478 418102
rect 565534 418046 565602 418102
rect 565658 418046 589194 418102
rect 589250 418046 589318 418102
rect 589374 418046 589442 418102
rect 589498 418046 589566 418102
rect 589622 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597980 418102
rect -1916 417978 597980 418046
rect -1916 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 5514 417978
rect 5570 417922 5638 417978
rect 5694 417922 5762 417978
rect 5818 417922 5886 417978
rect 5942 417922 12518 417978
rect 12574 417922 12642 417978
rect 12698 417922 43238 417978
rect 43294 417922 43362 417978
rect 43418 417922 73958 417978
rect 74014 417922 74082 417978
rect 74138 417922 104678 417978
rect 104734 417922 104802 417978
rect 104858 417922 135398 417978
rect 135454 417922 135522 417978
rect 135578 417922 166118 417978
rect 166174 417922 166242 417978
rect 166298 417922 196838 417978
rect 196894 417922 196962 417978
rect 197018 417922 227558 417978
rect 227614 417922 227682 417978
rect 227738 417922 258278 417978
rect 258334 417922 258402 417978
rect 258458 417922 288998 417978
rect 289054 417922 289122 417978
rect 289178 417922 319718 417978
rect 319774 417922 319842 417978
rect 319898 417922 350438 417978
rect 350494 417922 350562 417978
rect 350618 417922 381158 417978
rect 381214 417922 381282 417978
rect 381338 417922 411878 417978
rect 411934 417922 412002 417978
rect 412058 417922 442598 417978
rect 442654 417922 442722 417978
rect 442778 417922 473318 417978
rect 473374 417922 473442 417978
rect 473498 417922 504038 417978
rect 504094 417922 504162 417978
rect 504218 417922 534758 417978
rect 534814 417922 534882 417978
rect 534938 417922 565478 417978
rect 565534 417922 565602 417978
rect 565658 417922 589194 417978
rect 589250 417922 589318 417978
rect 589374 417922 589442 417978
rect 589498 417922 589566 417978
rect 589622 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597980 417978
rect -1916 417826 597980 417922
rect -1916 406350 597980 406446
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 27878 406350
rect 27934 406294 28002 406350
rect 28058 406294 58598 406350
rect 58654 406294 58722 406350
rect 58778 406294 89318 406350
rect 89374 406294 89442 406350
rect 89498 406294 120038 406350
rect 120094 406294 120162 406350
rect 120218 406294 150758 406350
rect 150814 406294 150882 406350
rect 150938 406294 181478 406350
rect 181534 406294 181602 406350
rect 181658 406294 212198 406350
rect 212254 406294 212322 406350
rect 212378 406294 242918 406350
rect 242974 406294 243042 406350
rect 243098 406294 273638 406350
rect 273694 406294 273762 406350
rect 273818 406294 304358 406350
rect 304414 406294 304482 406350
rect 304538 406294 335078 406350
rect 335134 406294 335202 406350
rect 335258 406294 365798 406350
rect 365854 406294 365922 406350
rect 365978 406294 396518 406350
rect 396574 406294 396642 406350
rect 396698 406294 427238 406350
rect 427294 406294 427362 406350
rect 427418 406294 457958 406350
rect 458014 406294 458082 406350
rect 458138 406294 488678 406350
rect 488734 406294 488802 406350
rect 488858 406294 519398 406350
rect 519454 406294 519522 406350
rect 519578 406294 550118 406350
rect 550174 406294 550242 406350
rect 550298 406294 592914 406350
rect 592970 406294 593038 406350
rect 593094 406294 593162 406350
rect 593218 406294 593286 406350
rect 593342 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect -1916 406226 597980 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 27878 406226
rect 27934 406170 28002 406226
rect 28058 406170 58598 406226
rect 58654 406170 58722 406226
rect 58778 406170 89318 406226
rect 89374 406170 89442 406226
rect 89498 406170 120038 406226
rect 120094 406170 120162 406226
rect 120218 406170 150758 406226
rect 150814 406170 150882 406226
rect 150938 406170 181478 406226
rect 181534 406170 181602 406226
rect 181658 406170 212198 406226
rect 212254 406170 212322 406226
rect 212378 406170 242918 406226
rect 242974 406170 243042 406226
rect 243098 406170 273638 406226
rect 273694 406170 273762 406226
rect 273818 406170 304358 406226
rect 304414 406170 304482 406226
rect 304538 406170 335078 406226
rect 335134 406170 335202 406226
rect 335258 406170 365798 406226
rect 365854 406170 365922 406226
rect 365978 406170 396518 406226
rect 396574 406170 396642 406226
rect 396698 406170 427238 406226
rect 427294 406170 427362 406226
rect 427418 406170 457958 406226
rect 458014 406170 458082 406226
rect 458138 406170 488678 406226
rect 488734 406170 488802 406226
rect 488858 406170 519398 406226
rect 519454 406170 519522 406226
rect 519578 406170 550118 406226
rect 550174 406170 550242 406226
rect 550298 406170 592914 406226
rect 592970 406170 593038 406226
rect 593094 406170 593162 406226
rect 593218 406170 593286 406226
rect 593342 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect -1916 406102 597980 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 27878 406102
rect 27934 406046 28002 406102
rect 28058 406046 58598 406102
rect 58654 406046 58722 406102
rect 58778 406046 89318 406102
rect 89374 406046 89442 406102
rect 89498 406046 120038 406102
rect 120094 406046 120162 406102
rect 120218 406046 150758 406102
rect 150814 406046 150882 406102
rect 150938 406046 181478 406102
rect 181534 406046 181602 406102
rect 181658 406046 212198 406102
rect 212254 406046 212322 406102
rect 212378 406046 242918 406102
rect 242974 406046 243042 406102
rect 243098 406046 273638 406102
rect 273694 406046 273762 406102
rect 273818 406046 304358 406102
rect 304414 406046 304482 406102
rect 304538 406046 335078 406102
rect 335134 406046 335202 406102
rect 335258 406046 365798 406102
rect 365854 406046 365922 406102
rect 365978 406046 396518 406102
rect 396574 406046 396642 406102
rect 396698 406046 427238 406102
rect 427294 406046 427362 406102
rect 427418 406046 457958 406102
rect 458014 406046 458082 406102
rect 458138 406046 488678 406102
rect 488734 406046 488802 406102
rect 488858 406046 519398 406102
rect 519454 406046 519522 406102
rect 519578 406046 550118 406102
rect 550174 406046 550242 406102
rect 550298 406046 592914 406102
rect 592970 406046 593038 406102
rect 593094 406046 593162 406102
rect 593218 406046 593286 406102
rect 593342 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect -1916 405978 597980 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 27878 405978
rect 27934 405922 28002 405978
rect 28058 405922 58598 405978
rect 58654 405922 58722 405978
rect 58778 405922 89318 405978
rect 89374 405922 89442 405978
rect 89498 405922 120038 405978
rect 120094 405922 120162 405978
rect 120218 405922 150758 405978
rect 150814 405922 150882 405978
rect 150938 405922 181478 405978
rect 181534 405922 181602 405978
rect 181658 405922 212198 405978
rect 212254 405922 212322 405978
rect 212378 405922 242918 405978
rect 242974 405922 243042 405978
rect 243098 405922 273638 405978
rect 273694 405922 273762 405978
rect 273818 405922 304358 405978
rect 304414 405922 304482 405978
rect 304538 405922 335078 405978
rect 335134 405922 335202 405978
rect 335258 405922 365798 405978
rect 365854 405922 365922 405978
rect 365978 405922 396518 405978
rect 396574 405922 396642 405978
rect 396698 405922 427238 405978
rect 427294 405922 427362 405978
rect 427418 405922 457958 405978
rect 458014 405922 458082 405978
rect 458138 405922 488678 405978
rect 488734 405922 488802 405978
rect 488858 405922 519398 405978
rect 519454 405922 519522 405978
rect 519578 405922 550118 405978
rect 550174 405922 550242 405978
rect 550298 405922 592914 405978
rect 592970 405922 593038 405978
rect 593094 405922 593162 405978
rect 593218 405922 593286 405978
rect 593342 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect -1916 405826 597980 405922
rect -1916 400350 597980 400446
rect -1916 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 5514 400350
rect 5570 400294 5638 400350
rect 5694 400294 5762 400350
rect 5818 400294 5886 400350
rect 5942 400294 12518 400350
rect 12574 400294 12642 400350
rect 12698 400294 43238 400350
rect 43294 400294 43362 400350
rect 43418 400294 73958 400350
rect 74014 400294 74082 400350
rect 74138 400294 104678 400350
rect 104734 400294 104802 400350
rect 104858 400294 135398 400350
rect 135454 400294 135522 400350
rect 135578 400294 166118 400350
rect 166174 400294 166242 400350
rect 166298 400294 196838 400350
rect 196894 400294 196962 400350
rect 197018 400294 227558 400350
rect 227614 400294 227682 400350
rect 227738 400294 258278 400350
rect 258334 400294 258402 400350
rect 258458 400294 288998 400350
rect 289054 400294 289122 400350
rect 289178 400294 319718 400350
rect 319774 400294 319842 400350
rect 319898 400294 350438 400350
rect 350494 400294 350562 400350
rect 350618 400294 381158 400350
rect 381214 400294 381282 400350
rect 381338 400294 411878 400350
rect 411934 400294 412002 400350
rect 412058 400294 442598 400350
rect 442654 400294 442722 400350
rect 442778 400294 473318 400350
rect 473374 400294 473442 400350
rect 473498 400294 504038 400350
rect 504094 400294 504162 400350
rect 504218 400294 534758 400350
rect 534814 400294 534882 400350
rect 534938 400294 565478 400350
rect 565534 400294 565602 400350
rect 565658 400294 589194 400350
rect 589250 400294 589318 400350
rect 589374 400294 589442 400350
rect 589498 400294 589566 400350
rect 589622 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597980 400350
rect -1916 400226 597980 400294
rect -1916 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 5514 400226
rect 5570 400170 5638 400226
rect 5694 400170 5762 400226
rect 5818 400170 5886 400226
rect 5942 400170 12518 400226
rect 12574 400170 12642 400226
rect 12698 400170 43238 400226
rect 43294 400170 43362 400226
rect 43418 400170 73958 400226
rect 74014 400170 74082 400226
rect 74138 400170 104678 400226
rect 104734 400170 104802 400226
rect 104858 400170 135398 400226
rect 135454 400170 135522 400226
rect 135578 400170 166118 400226
rect 166174 400170 166242 400226
rect 166298 400170 196838 400226
rect 196894 400170 196962 400226
rect 197018 400170 227558 400226
rect 227614 400170 227682 400226
rect 227738 400170 258278 400226
rect 258334 400170 258402 400226
rect 258458 400170 288998 400226
rect 289054 400170 289122 400226
rect 289178 400170 319718 400226
rect 319774 400170 319842 400226
rect 319898 400170 350438 400226
rect 350494 400170 350562 400226
rect 350618 400170 381158 400226
rect 381214 400170 381282 400226
rect 381338 400170 411878 400226
rect 411934 400170 412002 400226
rect 412058 400170 442598 400226
rect 442654 400170 442722 400226
rect 442778 400170 473318 400226
rect 473374 400170 473442 400226
rect 473498 400170 504038 400226
rect 504094 400170 504162 400226
rect 504218 400170 534758 400226
rect 534814 400170 534882 400226
rect 534938 400170 565478 400226
rect 565534 400170 565602 400226
rect 565658 400170 589194 400226
rect 589250 400170 589318 400226
rect 589374 400170 589442 400226
rect 589498 400170 589566 400226
rect 589622 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597980 400226
rect -1916 400102 597980 400170
rect -1916 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 5514 400102
rect 5570 400046 5638 400102
rect 5694 400046 5762 400102
rect 5818 400046 5886 400102
rect 5942 400046 12518 400102
rect 12574 400046 12642 400102
rect 12698 400046 43238 400102
rect 43294 400046 43362 400102
rect 43418 400046 73958 400102
rect 74014 400046 74082 400102
rect 74138 400046 104678 400102
rect 104734 400046 104802 400102
rect 104858 400046 135398 400102
rect 135454 400046 135522 400102
rect 135578 400046 166118 400102
rect 166174 400046 166242 400102
rect 166298 400046 196838 400102
rect 196894 400046 196962 400102
rect 197018 400046 227558 400102
rect 227614 400046 227682 400102
rect 227738 400046 258278 400102
rect 258334 400046 258402 400102
rect 258458 400046 288998 400102
rect 289054 400046 289122 400102
rect 289178 400046 319718 400102
rect 319774 400046 319842 400102
rect 319898 400046 350438 400102
rect 350494 400046 350562 400102
rect 350618 400046 381158 400102
rect 381214 400046 381282 400102
rect 381338 400046 411878 400102
rect 411934 400046 412002 400102
rect 412058 400046 442598 400102
rect 442654 400046 442722 400102
rect 442778 400046 473318 400102
rect 473374 400046 473442 400102
rect 473498 400046 504038 400102
rect 504094 400046 504162 400102
rect 504218 400046 534758 400102
rect 534814 400046 534882 400102
rect 534938 400046 565478 400102
rect 565534 400046 565602 400102
rect 565658 400046 589194 400102
rect 589250 400046 589318 400102
rect 589374 400046 589442 400102
rect 589498 400046 589566 400102
rect 589622 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597980 400102
rect -1916 399978 597980 400046
rect -1916 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 5514 399978
rect 5570 399922 5638 399978
rect 5694 399922 5762 399978
rect 5818 399922 5886 399978
rect 5942 399922 12518 399978
rect 12574 399922 12642 399978
rect 12698 399922 43238 399978
rect 43294 399922 43362 399978
rect 43418 399922 73958 399978
rect 74014 399922 74082 399978
rect 74138 399922 104678 399978
rect 104734 399922 104802 399978
rect 104858 399922 135398 399978
rect 135454 399922 135522 399978
rect 135578 399922 166118 399978
rect 166174 399922 166242 399978
rect 166298 399922 196838 399978
rect 196894 399922 196962 399978
rect 197018 399922 227558 399978
rect 227614 399922 227682 399978
rect 227738 399922 258278 399978
rect 258334 399922 258402 399978
rect 258458 399922 288998 399978
rect 289054 399922 289122 399978
rect 289178 399922 319718 399978
rect 319774 399922 319842 399978
rect 319898 399922 350438 399978
rect 350494 399922 350562 399978
rect 350618 399922 381158 399978
rect 381214 399922 381282 399978
rect 381338 399922 411878 399978
rect 411934 399922 412002 399978
rect 412058 399922 442598 399978
rect 442654 399922 442722 399978
rect 442778 399922 473318 399978
rect 473374 399922 473442 399978
rect 473498 399922 504038 399978
rect 504094 399922 504162 399978
rect 504218 399922 534758 399978
rect 534814 399922 534882 399978
rect 534938 399922 565478 399978
rect 565534 399922 565602 399978
rect 565658 399922 589194 399978
rect 589250 399922 589318 399978
rect 589374 399922 589442 399978
rect 589498 399922 589566 399978
rect 589622 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597980 399978
rect -1916 399826 597980 399922
rect -1916 388350 597980 388446
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 27878 388350
rect 27934 388294 28002 388350
rect 28058 388294 58598 388350
rect 58654 388294 58722 388350
rect 58778 388294 89318 388350
rect 89374 388294 89442 388350
rect 89498 388294 120038 388350
rect 120094 388294 120162 388350
rect 120218 388294 150758 388350
rect 150814 388294 150882 388350
rect 150938 388294 181478 388350
rect 181534 388294 181602 388350
rect 181658 388294 212198 388350
rect 212254 388294 212322 388350
rect 212378 388294 242918 388350
rect 242974 388294 243042 388350
rect 243098 388294 273638 388350
rect 273694 388294 273762 388350
rect 273818 388294 304358 388350
rect 304414 388294 304482 388350
rect 304538 388294 335078 388350
rect 335134 388294 335202 388350
rect 335258 388294 365798 388350
rect 365854 388294 365922 388350
rect 365978 388294 396518 388350
rect 396574 388294 396642 388350
rect 396698 388294 427238 388350
rect 427294 388294 427362 388350
rect 427418 388294 457958 388350
rect 458014 388294 458082 388350
rect 458138 388294 488678 388350
rect 488734 388294 488802 388350
rect 488858 388294 519398 388350
rect 519454 388294 519522 388350
rect 519578 388294 550118 388350
rect 550174 388294 550242 388350
rect 550298 388294 592914 388350
rect 592970 388294 593038 388350
rect 593094 388294 593162 388350
rect 593218 388294 593286 388350
rect 593342 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect -1916 388226 597980 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 27878 388226
rect 27934 388170 28002 388226
rect 28058 388170 58598 388226
rect 58654 388170 58722 388226
rect 58778 388170 89318 388226
rect 89374 388170 89442 388226
rect 89498 388170 120038 388226
rect 120094 388170 120162 388226
rect 120218 388170 150758 388226
rect 150814 388170 150882 388226
rect 150938 388170 181478 388226
rect 181534 388170 181602 388226
rect 181658 388170 212198 388226
rect 212254 388170 212322 388226
rect 212378 388170 242918 388226
rect 242974 388170 243042 388226
rect 243098 388170 273638 388226
rect 273694 388170 273762 388226
rect 273818 388170 304358 388226
rect 304414 388170 304482 388226
rect 304538 388170 335078 388226
rect 335134 388170 335202 388226
rect 335258 388170 365798 388226
rect 365854 388170 365922 388226
rect 365978 388170 396518 388226
rect 396574 388170 396642 388226
rect 396698 388170 427238 388226
rect 427294 388170 427362 388226
rect 427418 388170 457958 388226
rect 458014 388170 458082 388226
rect 458138 388170 488678 388226
rect 488734 388170 488802 388226
rect 488858 388170 519398 388226
rect 519454 388170 519522 388226
rect 519578 388170 550118 388226
rect 550174 388170 550242 388226
rect 550298 388170 592914 388226
rect 592970 388170 593038 388226
rect 593094 388170 593162 388226
rect 593218 388170 593286 388226
rect 593342 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect -1916 388102 597980 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 27878 388102
rect 27934 388046 28002 388102
rect 28058 388046 58598 388102
rect 58654 388046 58722 388102
rect 58778 388046 89318 388102
rect 89374 388046 89442 388102
rect 89498 388046 120038 388102
rect 120094 388046 120162 388102
rect 120218 388046 150758 388102
rect 150814 388046 150882 388102
rect 150938 388046 181478 388102
rect 181534 388046 181602 388102
rect 181658 388046 212198 388102
rect 212254 388046 212322 388102
rect 212378 388046 242918 388102
rect 242974 388046 243042 388102
rect 243098 388046 273638 388102
rect 273694 388046 273762 388102
rect 273818 388046 304358 388102
rect 304414 388046 304482 388102
rect 304538 388046 335078 388102
rect 335134 388046 335202 388102
rect 335258 388046 365798 388102
rect 365854 388046 365922 388102
rect 365978 388046 396518 388102
rect 396574 388046 396642 388102
rect 396698 388046 427238 388102
rect 427294 388046 427362 388102
rect 427418 388046 457958 388102
rect 458014 388046 458082 388102
rect 458138 388046 488678 388102
rect 488734 388046 488802 388102
rect 488858 388046 519398 388102
rect 519454 388046 519522 388102
rect 519578 388046 550118 388102
rect 550174 388046 550242 388102
rect 550298 388046 592914 388102
rect 592970 388046 593038 388102
rect 593094 388046 593162 388102
rect 593218 388046 593286 388102
rect 593342 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect -1916 387978 597980 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 27878 387978
rect 27934 387922 28002 387978
rect 28058 387922 58598 387978
rect 58654 387922 58722 387978
rect 58778 387922 89318 387978
rect 89374 387922 89442 387978
rect 89498 387922 120038 387978
rect 120094 387922 120162 387978
rect 120218 387922 150758 387978
rect 150814 387922 150882 387978
rect 150938 387922 181478 387978
rect 181534 387922 181602 387978
rect 181658 387922 212198 387978
rect 212254 387922 212322 387978
rect 212378 387922 242918 387978
rect 242974 387922 243042 387978
rect 243098 387922 273638 387978
rect 273694 387922 273762 387978
rect 273818 387922 304358 387978
rect 304414 387922 304482 387978
rect 304538 387922 335078 387978
rect 335134 387922 335202 387978
rect 335258 387922 365798 387978
rect 365854 387922 365922 387978
rect 365978 387922 396518 387978
rect 396574 387922 396642 387978
rect 396698 387922 427238 387978
rect 427294 387922 427362 387978
rect 427418 387922 457958 387978
rect 458014 387922 458082 387978
rect 458138 387922 488678 387978
rect 488734 387922 488802 387978
rect 488858 387922 519398 387978
rect 519454 387922 519522 387978
rect 519578 387922 550118 387978
rect 550174 387922 550242 387978
rect 550298 387922 592914 387978
rect 592970 387922 593038 387978
rect 593094 387922 593162 387978
rect 593218 387922 593286 387978
rect 593342 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect -1916 387826 597980 387922
rect -1916 382350 597980 382446
rect -1916 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 5514 382350
rect 5570 382294 5638 382350
rect 5694 382294 5762 382350
rect 5818 382294 5886 382350
rect 5942 382294 12518 382350
rect 12574 382294 12642 382350
rect 12698 382294 43238 382350
rect 43294 382294 43362 382350
rect 43418 382294 73958 382350
rect 74014 382294 74082 382350
rect 74138 382294 104678 382350
rect 104734 382294 104802 382350
rect 104858 382294 135398 382350
rect 135454 382294 135522 382350
rect 135578 382294 166118 382350
rect 166174 382294 166242 382350
rect 166298 382294 196838 382350
rect 196894 382294 196962 382350
rect 197018 382294 227558 382350
rect 227614 382294 227682 382350
rect 227738 382294 258278 382350
rect 258334 382294 258402 382350
rect 258458 382294 288998 382350
rect 289054 382294 289122 382350
rect 289178 382294 319718 382350
rect 319774 382294 319842 382350
rect 319898 382294 350438 382350
rect 350494 382294 350562 382350
rect 350618 382294 381158 382350
rect 381214 382294 381282 382350
rect 381338 382294 411878 382350
rect 411934 382294 412002 382350
rect 412058 382294 442598 382350
rect 442654 382294 442722 382350
rect 442778 382294 473318 382350
rect 473374 382294 473442 382350
rect 473498 382294 504038 382350
rect 504094 382294 504162 382350
rect 504218 382294 534758 382350
rect 534814 382294 534882 382350
rect 534938 382294 565478 382350
rect 565534 382294 565602 382350
rect 565658 382294 589194 382350
rect 589250 382294 589318 382350
rect 589374 382294 589442 382350
rect 589498 382294 589566 382350
rect 589622 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597980 382350
rect -1916 382226 597980 382294
rect -1916 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 5514 382226
rect 5570 382170 5638 382226
rect 5694 382170 5762 382226
rect 5818 382170 5886 382226
rect 5942 382170 12518 382226
rect 12574 382170 12642 382226
rect 12698 382170 43238 382226
rect 43294 382170 43362 382226
rect 43418 382170 73958 382226
rect 74014 382170 74082 382226
rect 74138 382170 104678 382226
rect 104734 382170 104802 382226
rect 104858 382170 135398 382226
rect 135454 382170 135522 382226
rect 135578 382170 166118 382226
rect 166174 382170 166242 382226
rect 166298 382170 196838 382226
rect 196894 382170 196962 382226
rect 197018 382170 227558 382226
rect 227614 382170 227682 382226
rect 227738 382170 258278 382226
rect 258334 382170 258402 382226
rect 258458 382170 288998 382226
rect 289054 382170 289122 382226
rect 289178 382170 319718 382226
rect 319774 382170 319842 382226
rect 319898 382170 350438 382226
rect 350494 382170 350562 382226
rect 350618 382170 381158 382226
rect 381214 382170 381282 382226
rect 381338 382170 411878 382226
rect 411934 382170 412002 382226
rect 412058 382170 442598 382226
rect 442654 382170 442722 382226
rect 442778 382170 473318 382226
rect 473374 382170 473442 382226
rect 473498 382170 504038 382226
rect 504094 382170 504162 382226
rect 504218 382170 534758 382226
rect 534814 382170 534882 382226
rect 534938 382170 565478 382226
rect 565534 382170 565602 382226
rect 565658 382170 589194 382226
rect 589250 382170 589318 382226
rect 589374 382170 589442 382226
rect 589498 382170 589566 382226
rect 589622 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597980 382226
rect -1916 382102 597980 382170
rect -1916 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 5514 382102
rect 5570 382046 5638 382102
rect 5694 382046 5762 382102
rect 5818 382046 5886 382102
rect 5942 382046 12518 382102
rect 12574 382046 12642 382102
rect 12698 382046 43238 382102
rect 43294 382046 43362 382102
rect 43418 382046 73958 382102
rect 74014 382046 74082 382102
rect 74138 382046 104678 382102
rect 104734 382046 104802 382102
rect 104858 382046 135398 382102
rect 135454 382046 135522 382102
rect 135578 382046 166118 382102
rect 166174 382046 166242 382102
rect 166298 382046 196838 382102
rect 196894 382046 196962 382102
rect 197018 382046 227558 382102
rect 227614 382046 227682 382102
rect 227738 382046 258278 382102
rect 258334 382046 258402 382102
rect 258458 382046 288998 382102
rect 289054 382046 289122 382102
rect 289178 382046 319718 382102
rect 319774 382046 319842 382102
rect 319898 382046 350438 382102
rect 350494 382046 350562 382102
rect 350618 382046 381158 382102
rect 381214 382046 381282 382102
rect 381338 382046 411878 382102
rect 411934 382046 412002 382102
rect 412058 382046 442598 382102
rect 442654 382046 442722 382102
rect 442778 382046 473318 382102
rect 473374 382046 473442 382102
rect 473498 382046 504038 382102
rect 504094 382046 504162 382102
rect 504218 382046 534758 382102
rect 534814 382046 534882 382102
rect 534938 382046 565478 382102
rect 565534 382046 565602 382102
rect 565658 382046 589194 382102
rect 589250 382046 589318 382102
rect 589374 382046 589442 382102
rect 589498 382046 589566 382102
rect 589622 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597980 382102
rect -1916 381978 597980 382046
rect -1916 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 5514 381978
rect 5570 381922 5638 381978
rect 5694 381922 5762 381978
rect 5818 381922 5886 381978
rect 5942 381922 12518 381978
rect 12574 381922 12642 381978
rect 12698 381922 43238 381978
rect 43294 381922 43362 381978
rect 43418 381922 73958 381978
rect 74014 381922 74082 381978
rect 74138 381922 104678 381978
rect 104734 381922 104802 381978
rect 104858 381922 135398 381978
rect 135454 381922 135522 381978
rect 135578 381922 166118 381978
rect 166174 381922 166242 381978
rect 166298 381922 196838 381978
rect 196894 381922 196962 381978
rect 197018 381922 227558 381978
rect 227614 381922 227682 381978
rect 227738 381922 258278 381978
rect 258334 381922 258402 381978
rect 258458 381922 288998 381978
rect 289054 381922 289122 381978
rect 289178 381922 319718 381978
rect 319774 381922 319842 381978
rect 319898 381922 350438 381978
rect 350494 381922 350562 381978
rect 350618 381922 381158 381978
rect 381214 381922 381282 381978
rect 381338 381922 411878 381978
rect 411934 381922 412002 381978
rect 412058 381922 442598 381978
rect 442654 381922 442722 381978
rect 442778 381922 473318 381978
rect 473374 381922 473442 381978
rect 473498 381922 504038 381978
rect 504094 381922 504162 381978
rect 504218 381922 534758 381978
rect 534814 381922 534882 381978
rect 534938 381922 565478 381978
rect 565534 381922 565602 381978
rect 565658 381922 589194 381978
rect 589250 381922 589318 381978
rect 589374 381922 589442 381978
rect 589498 381922 589566 381978
rect 589622 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597980 381978
rect -1916 381826 597980 381922
rect -1916 370350 597980 370446
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 27878 370350
rect 27934 370294 28002 370350
rect 28058 370294 58598 370350
rect 58654 370294 58722 370350
rect 58778 370294 89318 370350
rect 89374 370294 89442 370350
rect 89498 370294 120038 370350
rect 120094 370294 120162 370350
rect 120218 370294 150758 370350
rect 150814 370294 150882 370350
rect 150938 370294 181478 370350
rect 181534 370294 181602 370350
rect 181658 370294 212198 370350
rect 212254 370294 212322 370350
rect 212378 370294 242918 370350
rect 242974 370294 243042 370350
rect 243098 370294 273638 370350
rect 273694 370294 273762 370350
rect 273818 370294 304358 370350
rect 304414 370294 304482 370350
rect 304538 370294 335078 370350
rect 335134 370294 335202 370350
rect 335258 370294 365798 370350
rect 365854 370294 365922 370350
rect 365978 370294 396518 370350
rect 396574 370294 396642 370350
rect 396698 370294 427238 370350
rect 427294 370294 427362 370350
rect 427418 370294 457958 370350
rect 458014 370294 458082 370350
rect 458138 370294 488678 370350
rect 488734 370294 488802 370350
rect 488858 370294 519398 370350
rect 519454 370294 519522 370350
rect 519578 370294 550118 370350
rect 550174 370294 550242 370350
rect 550298 370294 592914 370350
rect 592970 370294 593038 370350
rect 593094 370294 593162 370350
rect 593218 370294 593286 370350
rect 593342 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect -1916 370226 597980 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 27878 370226
rect 27934 370170 28002 370226
rect 28058 370170 58598 370226
rect 58654 370170 58722 370226
rect 58778 370170 89318 370226
rect 89374 370170 89442 370226
rect 89498 370170 120038 370226
rect 120094 370170 120162 370226
rect 120218 370170 150758 370226
rect 150814 370170 150882 370226
rect 150938 370170 181478 370226
rect 181534 370170 181602 370226
rect 181658 370170 212198 370226
rect 212254 370170 212322 370226
rect 212378 370170 242918 370226
rect 242974 370170 243042 370226
rect 243098 370170 273638 370226
rect 273694 370170 273762 370226
rect 273818 370170 304358 370226
rect 304414 370170 304482 370226
rect 304538 370170 335078 370226
rect 335134 370170 335202 370226
rect 335258 370170 365798 370226
rect 365854 370170 365922 370226
rect 365978 370170 396518 370226
rect 396574 370170 396642 370226
rect 396698 370170 427238 370226
rect 427294 370170 427362 370226
rect 427418 370170 457958 370226
rect 458014 370170 458082 370226
rect 458138 370170 488678 370226
rect 488734 370170 488802 370226
rect 488858 370170 519398 370226
rect 519454 370170 519522 370226
rect 519578 370170 550118 370226
rect 550174 370170 550242 370226
rect 550298 370170 592914 370226
rect 592970 370170 593038 370226
rect 593094 370170 593162 370226
rect 593218 370170 593286 370226
rect 593342 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect -1916 370102 597980 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 27878 370102
rect 27934 370046 28002 370102
rect 28058 370046 58598 370102
rect 58654 370046 58722 370102
rect 58778 370046 89318 370102
rect 89374 370046 89442 370102
rect 89498 370046 120038 370102
rect 120094 370046 120162 370102
rect 120218 370046 150758 370102
rect 150814 370046 150882 370102
rect 150938 370046 181478 370102
rect 181534 370046 181602 370102
rect 181658 370046 212198 370102
rect 212254 370046 212322 370102
rect 212378 370046 242918 370102
rect 242974 370046 243042 370102
rect 243098 370046 273638 370102
rect 273694 370046 273762 370102
rect 273818 370046 304358 370102
rect 304414 370046 304482 370102
rect 304538 370046 335078 370102
rect 335134 370046 335202 370102
rect 335258 370046 365798 370102
rect 365854 370046 365922 370102
rect 365978 370046 396518 370102
rect 396574 370046 396642 370102
rect 396698 370046 427238 370102
rect 427294 370046 427362 370102
rect 427418 370046 457958 370102
rect 458014 370046 458082 370102
rect 458138 370046 488678 370102
rect 488734 370046 488802 370102
rect 488858 370046 519398 370102
rect 519454 370046 519522 370102
rect 519578 370046 550118 370102
rect 550174 370046 550242 370102
rect 550298 370046 592914 370102
rect 592970 370046 593038 370102
rect 593094 370046 593162 370102
rect 593218 370046 593286 370102
rect 593342 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect -1916 369978 597980 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 27878 369978
rect 27934 369922 28002 369978
rect 28058 369922 58598 369978
rect 58654 369922 58722 369978
rect 58778 369922 89318 369978
rect 89374 369922 89442 369978
rect 89498 369922 120038 369978
rect 120094 369922 120162 369978
rect 120218 369922 150758 369978
rect 150814 369922 150882 369978
rect 150938 369922 181478 369978
rect 181534 369922 181602 369978
rect 181658 369922 212198 369978
rect 212254 369922 212322 369978
rect 212378 369922 242918 369978
rect 242974 369922 243042 369978
rect 243098 369922 273638 369978
rect 273694 369922 273762 369978
rect 273818 369922 304358 369978
rect 304414 369922 304482 369978
rect 304538 369922 335078 369978
rect 335134 369922 335202 369978
rect 335258 369922 365798 369978
rect 365854 369922 365922 369978
rect 365978 369922 396518 369978
rect 396574 369922 396642 369978
rect 396698 369922 427238 369978
rect 427294 369922 427362 369978
rect 427418 369922 457958 369978
rect 458014 369922 458082 369978
rect 458138 369922 488678 369978
rect 488734 369922 488802 369978
rect 488858 369922 519398 369978
rect 519454 369922 519522 369978
rect 519578 369922 550118 369978
rect 550174 369922 550242 369978
rect 550298 369922 592914 369978
rect 592970 369922 593038 369978
rect 593094 369922 593162 369978
rect 593218 369922 593286 369978
rect 593342 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect -1916 369826 597980 369922
rect -1916 364350 597980 364446
rect -1916 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 5514 364350
rect 5570 364294 5638 364350
rect 5694 364294 5762 364350
rect 5818 364294 5886 364350
rect 5942 364294 12518 364350
rect 12574 364294 12642 364350
rect 12698 364294 43238 364350
rect 43294 364294 43362 364350
rect 43418 364294 73958 364350
rect 74014 364294 74082 364350
rect 74138 364294 104678 364350
rect 104734 364294 104802 364350
rect 104858 364294 135398 364350
rect 135454 364294 135522 364350
rect 135578 364294 166118 364350
rect 166174 364294 166242 364350
rect 166298 364294 196838 364350
rect 196894 364294 196962 364350
rect 197018 364294 227558 364350
rect 227614 364294 227682 364350
rect 227738 364294 258278 364350
rect 258334 364294 258402 364350
rect 258458 364294 288998 364350
rect 289054 364294 289122 364350
rect 289178 364294 319718 364350
rect 319774 364294 319842 364350
rect 319898 364294 350438 364350
rect 350494 364294 350562 364350
rect 350618 364294 381158 364350
rect 381214 364294 381282 364350
rect 381338 364294 411878 364350
rect 411934 364294 412002 364350
rect 412058 364294 442598 364350
rect 442654 364294 442722 364350
rect 442778 364294 473318 364350
rect 473374 364294 473442 364350
rect 473498 364294 504038 364350
rect 504094 364294 504162 364350
rect 504218 364294 534758 364350
rect 534814 364294 534882 364350
rect 534938 364294 565478 364350
rect 565534 364294 565602 364350
rect 565658 364294 589194 364350
rect 589250 364294 589318 364350
rect 589374 364294 589442 364350
rect 589498 364294 589566 364350
rect 589622 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597980 364350
rect -1916 364226 597980 364294
rect -1916 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 5514 364226
rect 5570 364170 5638 364226
rect 5694 364170 5762 364226
rect 5818 364170 5886 364226
rect 5942 364170 12518 364226
rect 12574 364170 12642 364226
rect 12698 364170 43238 364226
rect 43294 364170 43362 364226
rect 43418 364170 73958 364226
rect 74014 364170 74082 364226
rect 74138 364170 104678 364226
rect 104734 364170 104802 364226
rect 104858 364170 135398 364226
rect 135454 364170 135522 364226
rect 135578 364170 166118 364226
rect 166174 364170 166242 364226
rect 166298 364170 196838 364226
rect 196894 364170 196962 364226
rect 197018 364170 227558 364226
rect 227614 364170 227682 364226
rect 227738 364170 258278 364226
rect 258334 364170 258402 364226
rect 258458 364170 288998 364226
rect 289054 364170 289122 364226
rect 289178 364170 319718 364226
rect 319774 364170 319842 364226
rect 319898 364170 350438 364226
rect 350494 364170 350562 364226
rect 350618 364170 381158 364226
rect 381214 364170 381282 364226
rect 381338 364170 411878 364226
rect 411934 364170 412002 364226
rect 412058 364170 442598 364226
rect 442654 364170 442722 364226
rect 442778 364170 473318 364226
rect 473374 364170 473442 364226
rect 473498 364170 504038 364226
rect 504094 364170 504162 364226
rect 504218 364170 534758 364226
rect 534814 364170 534882 364226
rect 534938 364170 565478 364226
rect 565534 364170 565602 364226
rect 565658 364170 589194 364226
rect 589250 364170 589318 364226
rect 589374 364170 589442 364226
rect 589498 364170 589566 364226
rect 589622 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597980 364226
rect -1916 364102 597980 364170
rect -1916 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 5514 364102
rect 5570 364046 5638 364102
rect 5694 364046 5762 364102
rect 5818 364046 5886 364102
rect 5942 364046 12518 364102
rect 12574 364046 12642 364102
rect 12698 364046 43238 364102
rect 43294 364046 43362 364102
rect 43418 364046 73958 364102
rect 74014 364046 74082 364102
rect 74138 364046 104678 364102
rect 104734 364046 104802 364102
rect 104858 364046 135398 364102
rect 135454 364046 135522 364102
rect 135578 364046 166118 364102
rect 166174 364046 166242 364102
rect 166298 364046 196838 364102
rect 196894 364046 196962 364102
rect 197018 364046 227558 364102
rect 227614 364046 227682 364102
rect 227738 364046 258278 364102
rect 258334 364046 258402 364102
rect 258458 364046 288998 364102
rect 289054 364046 289122 364102
rect 289178 364046 319718 364102
rect 319774 364046 319842 364102
rect 319898 364046 350438 364102
rect 350494 364046 350562 364102
rect 350618 364046 381158 364102
rect 381214 364046 381282 364102
rect 381338 364046 411878 364102
rect 411934 364046 412002 364102
rect 412058 364046 442598 364102
rect 442654 364046 442722 364102
rect 442778 364046 473318 364102
rect 473374 364046 473442 364102
rect 473498 364046 504038 364102
rect 504094 364046 504162 364102
rect 504218 364046 534758 364102
rect 534814 364046 534882 364102
rect 534938 364046 565478 364102
rect 565534 364046 565602 364102
rect 565658 364046 589194 364102
rect 589250 364046 589318 364102
rect 589374 364046 589442 364102
rect 589498 364046 589566 364102
rect 589622 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597980 364102
rect -1916 363978 597980 364046
rect -1916 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 5514 363978
rect 5570 363922 5638 363978
rect 5694 363922 5762 363978
rect 5818 363922 5886 363978
rect 5942 363922 12518 363978
rect 12574 363922 12642 363978
rect 12698 363922 43238 363978
rect 43294 363922 43362 363978
rect 43418 363922 73958 363978
rect 74014 363922 74082 363978
rect 74138 363922 104678 363978
rect 104734 363922 104802 363978
rect 104858 363922 135398 363978
rect 135454 363922 135522 363978
rect 135578 363922 166118 363978
rect 166174 363922 166242 363978
rect 166298 363922 196838 363978
rect 196894 363922 196962 363978
rect 197018 363922 227558 363978
rect 227614 363922 227682 363978
rect 227738 363922 258278 363978
rect 258334 363922 258402 363978
rect 258458 363922 288998 363978
rect 289054 363922 289122 363978
rect 289178 363922 319718 363978
rect 319774 363922 319842 363978
rect 319898 363922 350438 363978
rect 350494 363922 350562 363978
rect 350618 363922 381158 363978
rect 381214 363922 381282 363978
rect 381338 363922 411878 363978
rect 411934 363922 412002 363978
rect 412058 363922 442598 363978
rect 442654 363922 442722 363978
rect 442778 363922 473318 363978
rect 473374 363922 473442 363978
rect 473498 363922 504038 363978
rect 504094 363922 504162 363978
rect 504218 363922 534758 363978
rect 534814 363922 534882 363978
rect 534938 363922 565478 363978
rect 565534 363922 565602 363978
rect 565658 363922 589194 363978
rect 589250 363922 589318 363978
rect 589374 363922 589442 363978
rect 589498 363922 589566 363978
rect 589622 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597980 363978
rect -1916 363826 597980 363922
rect -1916 352350 597980 352446
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 27878 352350
rect 27934 352294 28002 352350
rect 28058 352294 58598 352350
rect 58654 352294 58722 352350
rect 58778 352294 89318 352350
rect 89374 352294 89442 352350
rect 89498 352294 120038 352350
rect 120094 352294 120162 352350
rect 120218 352294 150758 352350
rect 150814 352294 150882 352350
rect 150938 352294 181478 352350
rect 181534 352294 181602 352350
rect 181658 352294 212198 352350
rect 212254 352294 212322 352350
rect 212378 352294 242918 352350
rect 242974 352294 243042 352350
rect 243098 352294 273638 352350
rect 273694 352294 273762 352350
rect 273818 352294 304358 352350
rect 304414 352294 304482 352350
rect 304538 352294 335078 352350
rect 335134 352294 335202 352350
rect 335258 352294 365798 352350
rect 365854 352294 365922 352350
rect 365978 352294 396518 352350
rect 396574 352294 396642 352350
rect 396698 352294 427238 352350
rect 427294 352294 427362 352350
rect 427418 352294 457958 352350
rect 458014 352294 458082 352350
rect 458138 352294 488678 352350
rect 488734 352294 488802 352350
rect 488858 352294 519398 352350
rect 519454 352294 519522 352350
rect 519578 352294 550118 352350
rect 550174 352294 550242 352350
rect 550298 352294 592914 352350
rect 592970 352294 593038 352350
rect 593094 352294 593162 352350
rect 593218 352294 593286 352350
rect 593342 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect -1916 352226 597980 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 27878 352226
rect 27934 352170 28002 352226
rect 28058 352170 58598 352226
rect 58654 352170 58722 352226
rect 58778 352170 89318 352226
rect 89374 352170 89442 352226
rect 89498 352170 120038 352226
rect 120094 352170 120162 352226
rect 120218 352170 150758 352226
rect 150814 352170 150882 352226
rect 150938 352170 181478 352226
rect 181534 352170 181602 352226
rect 181658 352170 212198 352226
rect 212254 352170 212322 352226
rect 212378 352170 242918 352226
rect 242974 352170 243042 352226
rect 243098 352170 273638 352226
rect 273694 352170 273762 352226
rect 273818 352170 304358 352226
rect 304414 352170 304482 352226
rect 304538 352170 335078 352226
rect 335134 352170 335202 352226
rect 335258 352170 365798 352226
rect 365854 352170 365922 352226
rect 365978 352170 396518 352226
rect 396574 352170 396642 352226
rect 396698 352170 427238 352226
rect 427294 352170 427362 352226
rect 427418 352170 457958 352226
rect 458014 352170 458082 352226
rect 458138 352170 488678 352226
rect 488734 352170 488802 352226
rect 488858 352170 519398 352226
rect 519454 352170 519522 352226
rect 519578 352170 550118 352226
rect 550174 352170 550242 352226
rect 550298 352170 592914 352226
rect 592970 352170 593038 352226
rect 593094 352170 593162 352226
rect 593218 352170 593286 352226
rect 593342 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect -1916 352102 597980 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 27878 352102
rect 27934 352046 28002 352102
rect 28058 352046 58598 352102
rect 58654 352046 58722 352102
rect 58778 352046 89318 352102
rect 89374 352046 89442 352102
rect 89498 352046 120038 352102
rect 120094 352046 120162 352102
rect 120218 352046 150758 352102
rect 150814 352046 150882 352102
rect 150938 352046 181478 352102
rect 181534 352046 181602 352102
rect 181658 352046 212198 352102
rect 212254 352046 212322 352102
rect 212378 352046 242918 352102
rect 242974 352046 243042 352102
rect 243098 352046 273638 352102
rect 273694 352046 273762 352102
rect 273818 352046 304358 352102
rect 304414 352046 304482 352102
rect 304538 352046 335078 352102
rect 335134 352046 335202 352102
rect 335258 352046 365798 352102
rect 365854 352046 365922 352102
rect 365978 352046 396518 352102
rect 396574 352046 396642 352102
rect 396698 352046 427238 352102
rect 427294 352046 427362 352102
rect 427418 352046 457958 352102
rect 458014 352046 458082 352102
rect 458138 352046 488678 352102
rect 488734 352046 488802 352102
rect 488858 352046 519398 352102
rect 519454 352046 519522 352102
rect 519578 352046 550118 352102
rect 550174 352046 550242 352102
rect 550298 352046 592914 352102
rect 592970 352046 593038 352102
rect 593094 352046 593162 352102
rect 593218 352046 593286 352102
rect 593342 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect -1916 351978 597980 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 27878 351978
rect 27934 351922 28002 351978
rect 28058 351922 58598 351978
rect 58654 351922 58722 351978
rect 58778 351922 89318 351978
rect 89374 351922 89442 351978
rect 89498 351922 120038 351978
rect 120094 351922 120162 351978
rect 120218 351922 150758 351978
rect 150814 351922 150882 351978
rect 150938 351922 181478 351978
rect 181534 351922 181602 351978
rect 181658 351922 212198 351978
rect 212254 351922 212322 351978
rect 212378 351922 242918 351978
rect 242974 351922 243042 351978
rect 243098 351922 273638 351978
rect 273694 351922 273762 351978
rect 273818 351922 304358 351978
rect 304414 351922 304482 351978
rect 304538 351922 335078 351978
rect 335134 351922 335202 351978
rect 335258 351922 365798 351978
rect 365854 351922 365922 351978
rect 365978 351922 396518 351978
rect 396574 351922 396642 351978
rect 396698 351922 427238 351978
rect 427294 351922 427362 351978
rect 427418 351922 457958 351978
rect 458014 351922 458082 351978
rect 458138 351922 488678 351978
rect 488734 351922 488802 351978
rect 488858 351922 519398 351978
rect 519454 351922 519522 351978
rect 519578 351922 550118 351978
rect 550174 351922 550242 351978
rect 550298 351922 592914 351978
rect 592970 351922 593038 351978
rect 593094 351922 593162 351978
rect 593218 351922 593286 351978
rect 593342 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect -1916 351826 597980 351922
rect -1916 346350 597980 346446
rect -1916 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 5514 346350
rect 5570 346294 5638 346350
rect 5694 346294 5762 346350
rect 5818 346294 5886 346350
rect 5942 346294 12518 346350
rect 12574 346294 12642 346350
rect 12698 346294 43238 346350
rect 43294 346294 43362 346350
rect 43418 346294 73958 346350
rect 74014 346294 74082 346350
rect 74138 346294 104678 346350
rect 104734 346294 104802 346350
rect 104858 346294 135398 346350
rect 135454 346294 135522 346350
rect 135578 346294 166118 346350
rect 166174 346294 166242 346350
rect 166298 346294 196838 346350
rect 196894 346294 196962 346350
rect 197018 346294 227558 346350
rect 227614 346294 227682 346350
rect 227738 346294 258278 346350
rect 258334 346294 258402 346350
rect 258458 346294 288998 346350
rect 289054 346294 289122 346350
rect 289178 346294 319718 346350
rect 319774 346294 319842 346350
rect 319898 346294 350438 346350
rect 350494 346294 350562 346350
rect 350618 346294 381158 346350
rect 381214 346294 381282 346350
rect 381338 346294 411878 346350
rect 411934 346294 412002 346350
rect 412058 346294 442598 346350
rect 442654 346294 442722 346350
rect 442778 346294 473318 346350
rect 473374 346294 473442 346350
rect 473498 346294 504038 346350
rect 504094 346294 504162 346350
rect 504218 346294 534758 346350
rect 534814 346294 534882 346350
rect 534938 346294 565478 346350
rect 565534 346294 565602 346350
rect 565658 346294 589194 346350
rect 589250 346294 589318 346350
rect 589374 346294 589442 346350
rect 589498 346294 589566 346350
rect 589622 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597980 346350
rect -1916 346226 597980 346294
rect -1916 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 5514 346226
rect 5570 346170 5638 346226
rect 5694 346170 5762 346226
rect 5818 346170 5886 346226
rect 5942 346170 12518 346226
rect 12574 346170 12642 346226
rect 12698 346170 43238 346226
rect 43294 346170 43362 346226
rect 43418 346170 73958 346226
rect 74014 346170 74082 346226
rect 74138 346170 104678 346226
rect 104734 346170 104802 346226
rect 104858 346170 135398 346226
rect 135454 346170 135522 346226
rect 135578 346170 166118 346226
rect 166174 346170 166242 346226
rect 166298 346170 196838 346226
rect 196894 346170 196962 346226
rect 197018 346170 227558 346226
rect 227614 346170 227682 346226
rect 227738 346170 258278 346226
rect 258334 346170 258402 346226
rect 258458 346170 288998 346226
rect 289054 346170 289122 346226
rect 289178 346170 319718 346226
rect 319774 346170 319842 346226
rect 319898 346170 350438 346226
rect 350494 346170 350562 346226
rect 350618 346170 381158 346226
rect 381214 346170 381282 346226
rect 381338 346170 411878 346226
rect 411934 346170 412002 346226
rect 412058 346170 442598 346226
rect 442654 346170 442722 346226
rect 442778 346170 473318 346226
rect 473374 346170 473442 346226
rect 473498 346170 504038 346226
rect 504094 346170 504162 346226
rect 504218 346170 534758 346226
rect 534814 346170 534882 346226
rect 534938 346170 565478 346226
rect 565534 346170 565602 346226
rect 565658 346170 589194 346226
rect 589250 346170 589318 346226
rect 589374 346170 589442 346226
rect 589498 346170 589566 346226
rect 589622 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597980 346226
rect -1916 346102 597980 346170
rect -1916 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 5514 346102
rect 5570 346046 5638 346102
rect 5694 346046 5762 346102
rect 5818 346046 5886 346102
rect 5942 346046 12518 346102
rect 12574 346046 12642 346102
rect 12698 346046 43238 346102
rect 43294 346046 43362 346102
rect 43418 346046 73958 346102
rect 74014 346046 74082 346102
rect 74138 346046 104678 346102
rect 104734 346046 104802 346102
rect 104858 346046 135398 346102
rect 135454 346046 135522 346102
rect 135578 346046 166118 346102
rect 166174 346046 166242 346102
rect 166298 346046 196838 346102
rect 196894 346046 196962 346102
rect 197018 346046 227558 346102
rect 227614 346046 227682 346102
rect 227738 346046 258278 346102
rect 258334 346046 258402 346102
rect 258458 346046 288998 346102
rect 289054 346046 289122 346102
rect 289178 346046 319718 346102
rect 319774 346046 319842 346102
rect 319898 346046 350438 346102
rect 350494 346046 350562 346102
rect 350618 346046 381158 346102
rect 381214 346046 381282 346102
rect 381338 346046 411878 346102
rect 411934 346046 412002 346102
rect 412058 346046 442598 346102
rect 442654 346046 442722 346102
rect 442778 346046 473318 346102
rect 473374 346046 473442 346102
rect 473498 346046 504038 346102
rect 504094 346046 504162 346102
rect 504218 346046 534758 346102
rect 534814 346046 534882 346102
rect 534938 346046 565478 346102
rect 565534 346046 565602 346102
rect 565658 346046 589194 346102
rect 589250 346046 589318 346102
rect 589374 346046 589442 346102
rect 589498 346046 589566 346102
rect 589622 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597980 346102
rect -1916 345978 597980 346046
rect -1916 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 5514 345978
rect 5570 345922 5638 345978
rect 5694 345922 5762 345978
rect 5818 345922 5886 345978
rect 5942 345922 12518 345978
rect 12574 345922 12642 345978
rect 12698 345922 43238 345978
rect 43294 345922 43362 345978
rect 43418 345922 73958 345978
rect 74014 345922 74082 345978
rect 74138 345922 104678 345978
rect 104734 345922 104802 345978
rect 104858 345922 135398 345978
rect 135454 345922 135522 345978
rect 135578 345922 166118 345978
rect 166174 345922 166242 345978
rect 166298 345922 196838 345978
rect 196894 345922 196962 345978
rect 197018 345922 227558 345978
rect 227614 345922 227682 345978
rect 227738 345922 258278 345978
rect 258334 345922 258402 345978
rect 258458 345922 288998 345978
rect 289054 345922 289122 345978
rect 289178 345922 319718 345978
rect 319774 345922 319842 345978
rect 319898 345922 350438 345978
rect 350494 345922 350562 345978
rect 350618 345922 381158 345978
rect 381214 345922 381282 345978
rect 381338 345922 411878 345978
rect 411934 345922 412002 345978
rect 412058 345922 442598 345978
rect 442654 345922 442722 345978
rect 442778 345922 473318 345978
rect 473374 345922 473442 345978
rect 473498 345922 504038 345978
rect 504094 345922 504162 345978
rect 504218 345922 534758 345978
rect 534814 345922 534882 345978
rect 534938 345922 565478 345978
rect 565534 345922 565602 345978
rect 565658 345922 589194 345978
rect 589250 345922 589318 345978
rect 589374 345922 589442 345978
rect 589498 345922 589566 345978
rect 589622 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597980 345978
rect -1916 345826 597980 345922
rect -1916 334350 597980 334446
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 27878 334350
rect 27934 334294 28002 334350
rect 28058 334294 58598 334350
rect 58654 334294 58722 334350
rect 58778 334294 89318 334350
rect 89374 334294 89442 334350
rect 89498 334294 120038 334350
rect 120094 334294 120162 334350
rect 120218 334294 150758 334350
rect 150814 334294 150882 334350
rect 150938 334294 181478 334350
rect 181534 334294 181602 334350
rect 181658 334294 212198 334350
rect 212254 334294 212322 334350
rect 212378 334294 242918 334350
rect 242974 334294 243042 334350
rect 243098 334294 273638 334350
rect 273694 334294 273762 334350
rect 273818 334294 304358 334350
rect 304414 334294 304482 334350
rect 304538 334294 335078 334350
rect 335134 334294 335202 334350
rect 335258 334294 365798 334350
rect 365854 334294 365922 334350
rect 365978 334294 396518 334350
rect 396574 334294 396642 334350
rect 396698 334294 427238 334350
rect 427294 334294 427362 334350
rect 427418 334294 457958 334350
rect 458014 334294 458082 334350
rect 458138 334294 488678 334350
rect 488734 334294 488802 334350
rect 488858 334294 519398 334350
rect 519454 334294 519522 334350
rect 519578 334294 550118 334350
rect 550174 334294 550242 334350
rect 550298 334294 592914 334350
rect 592970 334294 593038 334350
rect 593094 334294 593162 334350
rect 593218 334294 593286 334350
rect 593342 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect -1916 334226 597980 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 27878 334226
rect 27934 334170 28002 334226
rect 28058 334170 58598 334226
rect 58654 334170 58722 334226
rect 58778 334170 89318 334226
rect 89374 334170 89442 334226
rect 89498 334170 120038 334226
rect 120094 334170 120162 334226
rect 120218 334170 150758 334226
rect 150814 334170 150882 334226
rect 150938 334170 181478 334226
rect 181534 334170 181602 334226
rect 181658 334170 212198 334226
rect 212254 334170 212322 334226
rect 212378 334170 242918 334226
rect 242974 334170 243042 334226
rect 243098 334170 273638 334226
rect 273694 334170 273762 334226
rect 273818 334170 304358 334226
rect 304414 334170 304482 334226
rect 304538 334170 335078 334226
rect 335134 334170 335202 334226
rect 335258 334170 365798 334226
rect 365854 334170 365922 334226
rect 365978 334170 396518 334226
rect 396574 334170 396642 334226
rect 396698 334170 427238 334226
rect 427294 334170 427362 334226
rect 427418 334170 457958 334226
rect 458014 334170 458082 334226
rect 458138 334170 488678 334226
rect 488734 334170 488802 334226
rect 488858 334170 519398 334226
rect 519454 334170 519522 334226
rect 519578 334170 550118 334226
rect 550174 334170 550242 334226
rect 550298 334170 592914 334226
rect 592970 334170 593038 334226
rect 593094 334170 593162 334226
rect 593218 334170 593286 334226
rect 593342 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect -1916 334102 597980 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 27878 334102
rect 27934 334046 28002 334102
rect 28058 334046 58598 334102
rect 58654 334046 58722 334102
rect 58778 334046 89318 334102
rect 89374 334046 89442 334102
rect 89498 334046 120038 334102
rect 120094 334046 120162 334102
rect 120218 334046 150758 334102
rect 150814 334046 150882 334102
rect 150938 334046 181478 334102
rect 181534 334046 181602 334102
rect 181658 334046 212198 334102
rect 212254 334046 212322 334102
rect 212378 334046 242918 334102
rect 242974 334046 243042 334102
rect 243098 334046 273638 334102
rect 273694 334046 273762 334102
rect 273818 334046 304358 334102
rect 304414 334046 304482 334102
rect 304538 334046 335078 334102
rect 335134 334046 335202 334102
rect 335258 334046 365798 334102
rect 365854 334046 365922 334102
rect 365978 334046 396518 334102
rect 396574 334046 396642 334102
rect 396698 334046 427238 334102
rect 427294 334046 427362 334102
rect 427418 334046 457958 334102
rect 458014 334046 458082 334102
rect 458138 334046 488678 334102
rect 488734 334046 488802 334102
rect 488858 334046 519398 334102
rect 519454 334046 519522 334102
rect 519578 334046 550118 334102
rect 550174 334046 550242 334102
rect 550298 334046 592914 334102
rect 592970 334046 593038 334102
rect 593094 334046 593162 334102
rect 593218 334046 593286 334102
rect 593342 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect -1916 333978 597980 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 27878 333978
rect 27934 333922 28002 333978
rect 28058 333922 58598 333978
rect 58654 333922 58722 333978
rect 58778 333922 89318 333978
rect 89374 333922 89442 333978
rect 89498 333922 120038 333978
rect 120094 333922 120162 333978
rect 120218 333922 150758 333978
rect 150814 333922 150882 333978
rect 150938 333922 181478 333978
rect 181534 333922 181602 333978
rect 181658 333922 212198 333978
rect 212254 333922 212322 333978
rect 212378 333922 242918 333978
rect 242974 333922 243042 333978
rect 243098 333922 273638 333978
rect 273694 333922 273762 333978
rect 273818 333922 304358 333978
rect 304414 333922 304482 333978
rect 304538 333922 335078 333978
rect 335134 333922 335202 333978
rect 335258 333922 365798 333978
rect 365854 333922 365922 333978
rect 365978 333922 396518 333978
rect 396574 333922 396642 333978
rect 396698 333922 427238 333978
rect 427294 333922 427362 333978
rect 427418 333922 457958 333978
rect 458014 333922 458082 333978
rect 458138 333922 488678 333978
rect 488734 333922 488802 333978
rect 488858 333922 519398 333978
rect 519454 333922 519522 333978
rect 519578 333922 550118 333978
rect 550174 333922 550242 333978
rect 550298 333922 592914 333978
rect 592970 333922 593038 333978
rect 593094 333922 593162 333978
rect 593218 333922 593286 333978
rect 593342 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect -1916 333826 597980 333922
rect -1916 328350 597980 328446
rect -1916 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 5514 328350
rect 5570 328294 5638 328350
rect 5694 328294 5762 328350
rect 5818 328294 5886 328350
rect 5942 328294 12518 328350
rect 12574 328294 12642 328350
rect 12698 328294 43238 328350
rect 43294 328294 43362 328350
rect 43418 328294 73958 328350
rect 74014 328294 74082 328350
rect 74138 328294 104678 328350
rect 104734 328294 104802 328350
rect 104858 328294 135398 328350
rect 135454 328294 135522 328350
rect 135578 328294 166118 328350
rect 166174 328294 166242 328350
rect 166298 328294 196838 328350
rect 196894 328294 196962 328350
rect 197018 328294 227558 328350
rect 227614 328294 227682 328350
rect 227738 328294 258278 328350
rect 258334 328294 258402 328350
rect 258458 328294 288998 328350
rect 289054 328294 289122 328350
rect 289178 328294 319718 328350
rect 319774 328294 319842 328350
rect 319898 328294 350438 328350
rect 350494 328294 350562 328350
rect 350618 328294 381158 328350
rect 381214 328294 381282 328350
rect 381338 328294 411878 328350
rect 411934 328294 412002 328350
rect 412058 328294 442598 328350
rect 442654 328294 442722 328350
rect 442778 328294 473318 328350
rect 473374 328294 473442 328350
rect 473498 328294 504038 328350
rect 504094 328294 504162 328350
rect 504218 328294 534758 328350
rect 534814 328294 534882 328350
rect 534938 328294 565478 328350
rect 565534 328294 565602 328350
rect 565658 328294 589194 328350
rect 589250 328294 589318 328350
rect 589374 328294 589442 328350
rect 589498 328294 589566 328350
rect 589622 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597980 328350
rect -1916 328226 597980 328294
rect -1916 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 5514 328226
rect 5570 328170 5638 328226
rect 5694 328170 5762 328226
rect 5818 328170 5886 328226
rect 5942 328170 12518 328226
rect 12574 328170 12642 328226
rect 12698 328170 43238 328226
rect 43294 328170 43362 328226
rect 43418 328170 73958 328226
rect 74014 328170 74082 328226
rect 74138 328170 104678 328226
rect 104734 328170 104802 328226
rect 104858 328170 135398 328226
rect 135454 328170 135522 328226
rect 135578 328170 166118 328226
rect 166174 328170 166242 328226
rect 166298 328170 196838 328226
rect 196894 328170 196962 328226
rect 197018 328170 227558 328226
rect 227614 328170 227682 328226
rect 227738 328170 258278 328226
rect 258334 328170 258402 328226
rect 258458 328170 288998 328226
rect 289054 328170 289122 328226
rect 289178 328170 319718 328226
rect 319774 328170 319842 328226
rect 319898 328170 350438 328226
rect 350494 328170 350562 328226
rect 350618 328170 381158 328226
rect 381214 328170 381282 328226
rect 381338 328170 411878 328226
rect 411934 328170 412002 328226
rect 412058 328170 442598 328226
rect 442654 328170 442722 328226
rect 442778 328170 473318 328226
rect 473374 328170 473442 328226
rect 473498 328170 504038 328226
rect 504094 328170 504162 328226
rect 504218 328170 534758 328226
rect 534814 328170 534882 328226
rect 534938 328170 565478 328226
rect 565534 328170 565602 328226
rect 565658 328170 589194 328226
rect 589250 328170 589318 328226
rect 589374 328170 589442 328226
rect 589498 328170 589566 328226
rect 589622 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597980 328226
rect -1916 328102 597980 328170
rect -1916 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 5514 328102
rect 5570 328046 5638 328102
rect 5694 328046 5762 328102
rect 5818 328046 5886 328102
rect 5942 328046 12518 328102
rect 12574 328046 12642 328102
rect 12698 328046 43238 328102
rect 43294 328046 43362 328102
rect 43418 328046 73958 328102
rect 74014 328046 74082 328102
rect 74138 328046 104678 328102
rect 104734 328046 104802 328102
rect 104858 328046 135398 328102
rect 135454 328046 135522 328102
rect 135578 328046 166118 328102
rect 166174 328046 166242 328102
rect 166298 328046 196838 328102
rect 196894 328046 196962 328102
rect 197018 328046 227558 328102
rect 227614 328046 227682 328102
rect 227738 328046 258278 328102
rect 258334 328046 258402 328102
rect 258458 328046 288998 328102
rect 289054 328046 289122 328102
rect 289178 328046 319718 328102
rect 319774 328046 319842 328102
rect 319898 328046 350438 328102
rect 350494 328046 350562 328102
rect 350618 328046 381158 328102
rect 381214 328046 381282 328102
rect 381338 328046 411878 328102
rect 411934 328046 412002 328102
rect 412058 328046 442598 328102
rect 442654 328046 442722 328102
rect 442778 328046 473318 328102
rect 473374 328046 473442 328102
rect 473498 328046 504038 328102
rect 504094 328046 504162 328102
rect 504218 328046 534758 328102
rect 534814 328046 534882 328102
rect 534938 328046 565478 328102
rect 565534 328046 565602 328102
rect 565658 328046 589194 328102
rect 589250 328046 589318 328102
rect 589374 328046 589442 328102
rect 589498 328046 589566 328102
rect 589622 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597980 328102
rect -1916 327978 597980 328046
rect -1916 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 5514 327978
rect 5570 327922 5638 327978
rect 5694 327922 5762 327978
rect 5818 327922 5886 327978
rect 5942 327922 12518 327978
rect 12574 327922 12642 327978
rect 12698 327922 43238 327978
rect 43294 327922 43362 327978
rect 43418 327922 73958 327978
rect 74014 327922 74082 327978
rect 74138 327922 104678 327978
rect 104734 327922 104802 327978
rect 104858 327922 135398 327978
rect 135454 327922 135522 327978
rect 135578 327922 166118 327978
rect 166174 327922 166242 327978
rect 166298 327922 196838 327978
rect 196894 327922 196962 327978
rect 197018 327922 227558 327978
rect 227614 327922 227682 327978
rect 227738 327922 258278 327978
rect 258334 327922 258402 327978
rect 258458 327922 288998 327978
rect 289054 327922 289122 327978
rect 289178 327922 319718 327978
rect 319774 327922 319842 327978
rect 319898 327922 350438 327978
rect 350494 327922 350562 327978
rect 350618 327922 381158 327978
rect 381214 327922 381282 327978
rect 381338 327922 411878 327978
rect 411934 327922 412002 327978
rect 412058 327922 442598 327978
rect 442654 327922 442722 327978
rect 442778 327922 473318 327978
rect 473374 327922 473442 327978
rect 473498 327922 504038 327978
rect 504094 327922 504162 327978
rect 504218 327922 534758 327978
rect 534814 327922 534882 327978
rect 534938 327922 565478 327978
rect 565534 327922 565602 327978
rect 565658 327922 589194 327978
rect 589250 327922 589318 327978
rect 589374 327922 589442 327978
rect 589498 327922 589566 327978
rect 589622 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597980 327978
rect -1916 327826 597980 327922
rect -1916 316350 597980 316446
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 27878 316350
rect 27934 316294 28002 316350
rect 28058 316294 58598 316350
rect 58654 316294 58722 316350
rect 58778 316294 89318 316350
rect 89374 316294 89442 316350
rect 89498 316294 120038 316350
rect 120094 316294 120162 316350
rect 120218 316294 150758 316350
rect 150814 316294 150882 316350
rect 150938 316294 181478 316350
rect 181534 316294 181602 316350
rect 181658 316294 212198 316350
rect 212254 316294 212322 316350
rect 212378 316294 242918 316350
rect 242974 316294 243042 316350
rect 243098 316294 273638 316350
rect 273694 316294 273762 316350
rect 273818 316294 304358 316350
rect 304414 316294 304482 316350
rect 304538 316294 335078 316350
rect 335134 316294 335202 316350
rect 335258 316294 365798 316350
rect 365854 316294 365922 316350
rect 365978 316294 396518 316350
rect 396574 316294 396642 316350
rect 396698 316294 427238 316350
rect 427294 316294 427362 316350
rect 427418 316294 457958 316350
rect 458014 316294 458082 316350
rect 458138 316294 488678 316350
rect 488734 316294 488802 316350
rect 488858 316294 519398 316350
rect 519454 316294 519522 316350
rect 519578 316294 550118 316350
rect 550174 316294 550242 316350
rect 550298 316294 592914 316350
rect 592970 316294 593038 316350
rect 593094 316294 593162 316350
rect 593218 316294 593286 316350
rect 593342 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect -1916 316226 597980 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 27878 316226
rect 27934 316170 28002 316226
rect 28058 316170 58598 316226
rect 58654 316170 58722 316226
rect 58778 316170 89318 316226
rect 89374 316170 89442 316226
rect 89498 316170 120038 316226
rect 120094 316170 120162 316226
rect 120218 316170 150758 316226
rect 150814 316170 150882 316226
rect 150938 316170 181478 316226
rect 181534 316170 181602 316226
rect 181658 316170 212198 316226
rect 212254 316170 212322 316226
rect 212378 316170 242918 316226
rect 242974 316170 243042 316226
rect 243098 316170 273638 316226
rect 273694 316170 273762 316226
rect 273818 316170 304358 316226
rect 304414 316170 304482 316226
rect 304538 316170 335078 316226
rect 335134 316170 335202 316226
rect 335258 316170 365798 316226
rect 365854 316170 365922 316226
rect 365978 316170 396518 316226
rect 396574 316170 396642 316226
rect 396698 316170 427238 316226
rect 427294 316170 427362 316226
rect 427418 316170 457958 316226
rect 458014 316170 458082 316226
rect 458138 316170 488678 316226
rect 488734 316170 488802 316226
rect 488858 316170 519398 316226
rect 519454 316170 519522 316226
rect 519578 316170 550118 316226
rect 550174 316170 550242 316226
rect 550298 316170 592914 316226
rect 592970 316170 593038 316226
rect 593094 316170 593162 316226
rect 593218 316170 593286 316226
rect 593342 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect -1916 316102 597980 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 27878 316102
rect 27934 316046 28002 316102
rect 28058 316046 58598 316102
rect 58654 316046 58722 316102
rect 58778 316046 89318 316102
rect 89374 316046 89442 316102
rect 89498 316046 120038 316102
rect 120094 316046 120162 316102
rect 120218 316046 150758 316102
rect 150814 316046 150882 316102
rect 150938 316046 181478 316102
rect 181534 316046 181602 316102
rect 181658 316046 212198 316102
rect 212254 316046 212322 316102
rect 212378 316046 242918 316102
rect 242974 316046 243042 316102
rect 243098 316046 273638 316102
rect 273694 316046 273762 316102
rect 273818 316046 304358 316102
rect 304414 316046 304482 316102
rect 304538 316046 335078 316102
rect 335134 316046 335202 316102
rect 335258 316046 365798 316102
rect 365854 316046 365922 316102
rect 365978 316046 396518 316102
rect 396574 316046 396642 316102
rect 396698 316046 427238 316102
rect 427294 316046 427362 316102
rect 427418 316046 457958 316102
rect 458014 316046 458082 316102
rect 458138 316046 488678 316102
rect 488734 316046 488802 316102
rect 488858 316046 519398 316102
rect 519454 316046 519522 316102
rect 519578 316046 550118 316102
rect 550174 316046 550242 316102
rect 550298 316046 592914 316102
rect 592970 316046 593038 316102
rect 593094 316046 593162 316102
rect 593218 316046 593286 316102
rect 593342 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect -1916 315978 597980 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 27878 315978
rect 27934 315922 28002 315978
rect 28058 315922 58598 315978
rect 58654 315922 58722 315978
rect 58778 315922 89318 315978
rect 89374 315922 89442 315978
rect 89498 315922 120038 315978
rect 120094 315922 120162 315978
rect 120218 315922 150758 315978
rect 150814 315922 150882 315978
rect 150938 315922 181478 315978
rect 181534 315922 181602 315978
rect 181658 315922 212198 315978
rect 212254 315922 212322 315978
rect 212378 315922 242918 315978
rect 242974 315922 243042 315978
rect 243098 315922 273638 315978
rect 273694 315922 273762 315978
rect 273818 315922 304358 315978
rect 304414 315922 304482 315978
rect 304538 315922 335078 315978
rect 335134 315922 335202 315978
rect 335258 315922 365798 315978
rect 365854 315922 365922 315978
rect 365978 315922 396518 315978
rect 396574 315922 396642 315978
rect 396698 315922 427238 315978
rect 427294 315922 427362 315978
rect 427418 315922 457958 315978
rect 458014 315922 458082 315978
rect 458138 315922 488678 315978
rect 488734 315922 488802 315978
rect 488858 315922 519398 315978
rect 519454 315922 519522 315978
rect 519578 315922 550118 315978
rect 550174 315922 550242 315978
rect 550298 315922 592914 315978
rect 592970 315922 593038 315978
rect 593094 315922 593162 315978
rect 593218 315922 593286 315978
rect 593342 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect -1916 315826 597980 315922
rect -1916 310350 597980 310446
rect -1916 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 5514 310350
rect 5570 310294 5638 310350
rect 5694 310294 5762 310350
rect 5818 310294 5886 310350
rect 5942 310294 12518 310350
rect 12574 310294 12642 310350
rect 12698 310294 43238 310350
rect 43294 310294 43362 310350
rect 43418 310294 73958 310350
rect 74014 310294 74082 310350
rect 74138 310294 104678 310350
rect 104734 310294 104802 310350
rect 104858 310294 135398 310350
rect 135454 310294 135522 310350
rect 135578 310294 166118 310350
rect 166174 310294 166242 310350
rect 166298 310294 196838 310350
rect 196894 310294 196962 310350
rect 197018 310294 227558 310350
rect 227614 310294 227682 310350
rect 227738 310294 258278 310350
rect 258334 310294 258402 310350
rect 258458 310294 288998 310350
rect 289054 310294 289122 310350
rect 289178 310294 319718 310350
rect 319774 310294 319842 310350
rect 319898 310294 350438 310350
rect 350494 310294 350562 310350
rect 350618 310294 381158 310350
rect 381214 310294 381282 310350
rect 381338 310294 411878 310350
rect 411934 310294 412002 310350
rect 412058 310294 442598 310350
rect 442654 310294 442722 310350
rect 442778 310294 473318 310350
rect 473374 310294 473442 310350
rect 473498 310294 504038 310350
rect 504094 310294 504162 310350
rect 504218 310294 534758 310350
rect 534814 310294 534882 310350
rect 534938 310294 565478 310350
rect 565534 310294 565602 310350
rect 565658 310294 589194 310350
rect 589250 310294 589318 310350
rect 589374 310294 589442 310350
rect 589498 310294 589566 310350
rect 589622 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597980 310350
rect -1916 310226 597980 310294
rect -1916 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 5514 310226
rect 5570 310170 5638 310226
rect 5694 310170 5762 310226
rect 5818 310170 5886 310226
rect 5942 310170 12518 310226
rect 12574 310170 12642 310226
rect 12698 310170 43238 310226
rect 43294 310170 43362 310226
rect 43418 310170 73958 310226
rect 74014 310170 74082 310226
rect 74138 310170 104678 310226
rect 104734 310170 104802 310226
rect 104858 310170 135398 310226
rect 135454 310170 135522 310226
rect 135578 310170 166118 310226
rect 166174 310170 166242 310226
rect 166298 310170 196838 310226
rect 196894 310170 196962 310226
rect 197018 310170 227558 310226
rect 227614 310170 227682 310226
rect 227738 310170 258278 310226
rect 258334 310170 258402 310226
rect 258458 310170 288998 310226
rect 289054 310170 289122 310226
rect 289178 310170 319718 310226
rect 319774 310170 319842 310226
rect 319898 310170 350438 310226
rect 350494 310170 350562 310226
rect 350618 310170 381158 310226
rect 381214 310170 381282 310226
rect 381338 310170 411878 310226
rect 411934 310170 412002 310226
rect 412058 310170 442598 310226
rect 442654 310170 442722 310226
rect 442778 310170 473318 310226
rect 473374 310170 473442 310226
rect 473498 310170 504038 310226
rect 504094 310170 504162 310226
rect 504218 310170 534758 310226
rect 534814 310170 534882 310226
rect 534938 310170 565478 310226
rect 565534 310170 565602 310226
rect 565658 310170 589194 310226
rect 589250 310170 589318 310226
rect 589374 310170 589442 310226
rect 589498 310170 589566 310226
rect 589622 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597980 310226
rect -1916 310102 597980 310170
rect -1916 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 5514 310102
rect 5570 310046 5638 310102
rect 5694 310046 5762 310102
rect 5818 310046 5886 310102
rect 5942 310046 12518 310102
rect 12574 310046 12642 310102
rect 12698 310046 43238 310102
rect 43294 310046 43362 310102
rect 43418 310046 73958 310102
rect 74014 310046 74082 310102
rect 74138 310046 104678 310102
rect 104734 310046 104802 310102
rect 104858 310046 135398 310102
rect 135454 310046 135522 310102
rect 135578 310046 166118 310102
rect 166174 310046 166242 310102
rect 166298 310046 196838 310102
rect 196894 310046 196962 310102
rect 197018 310046 227558 310102
rect 227614 310046 227682 310102
rect 227738 310046 258278 310102
rect 258334 310046 258402 310102
rect 258458 310046 288998 310102
rect 289054 310046 289122 310102
rect 289178 310046 319718 310102
rect 319774 310046 319842 310102
rect 319898 310046 350438 310102
rect 350494 310046 350562 310102
rect 350618 310046 381158 310102
rect 381214 310046 381282 310102
rect 381338 310046 411878 310102
rect 411934 310046 412002 310102
rect 412058 310046 442598 310102
rect 442654 310046 442722 310102
rect 442778 310046 473318 310102
rect 473374 310046 473442 310102
rect 473498 310046 504038 310102
rect 504094 310046 504162 310102
rect 504218 310046 534758 310102
rect 534814 310046 534882 310102
rect 534938 310046 565478 310102
rect 565534 310046 565602 310102
rect 565658 310046 589194 310102
rect 589250 310046 589318 310102
rect 589374 310046 589442 310102
rect 589498 310046 589566 310102
rect 589622 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597980 310102
rect -1916 309978 597980 310046
rect -1916 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 5514 309978
rect 5570 309922 5638 309978
rect 5694 309922 5762 309978
rect 5818 309922 5886 309978
rect 5942 309922 12518 309978
rect 12574 309922 12642 309978
rect 12698 309922 43238 309978
rect 43294 309922 43362 309978
rect 43418 309922 73958 309978
rect 74014 309922 74082 309978
rect 74138 309922 104678 309978
rect 104734 309922 104802 309978
rect 104858 309922 135398 309978
rect 135454 309922 135522 309978
rect 135578 309922 166118 309978
rect 166174 309922 166242 309978
rect 166298 309922 196838 309978
rect 196894 309922 196962 309978
rect 197018 309922 227558 309978
rect 227614 309922 227682 309978
rect 227738 309922 258278 309978
rect 258334 309922 258402 309978
rect 258458 309922 288998 309978
rect 289054 309922 289122 309978
rect 289178 309922 319718 309978
rect 319774 309922 319842 309978
rect 319898 309922 350438 309978
rect 350494 309922 350562 309978
rect 350618 309922 381158 309978
rect 381214 309922 381282 309978
rect 381338 309922 411878 309978
rect 411934 309922 412002 309978
rect 412058 309922 442598 309978
rect 442654 309922 442722 309978
rect 442778 309922 473318 309978
rect 473374 309922 473442 309978
rect 473498 309922 504038 309978
rect 504094 309922 504162 309978
rect 504218 309922 534758 309978
rect 534814 309922 534882 309978
rect 534938 309922 565478 309978
rect 565534 309922 565602 309978
rect 565658 309922 589194 309978
rect 589250 309922 589318 309978
rect 589374 309922 589442 309978
rect 589498 309922 589566 309978
rect 589622 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597980 309978
rect -1916 309826 597980 309922
rect -1916 298350 597980 298446
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 27878 298350
rect 27934 298294 28002 298350
rect 28058 298294 58598 298350
rect 58654 298294 58722 298350
rect 58778 298294 89318 298350
rect 89374 298294 89442 298350
rect 89498 298294 120038 298350
rect 120094 298294 120162 298350
rect 120218 298294 150758 298350
rect 150814 298294 150882 298350
rect 150938 298294 181478 298350
rect 181534 298294 181602 298350
rect 181658 298294 212198 298350
rect 212254 298294 212322 298350
rect 212378 298294 242918 298350
rect 242974 298294 243042 298350
rect 243098 298294 273638 298350
rect 273694 298294 273762 298350
rect 273818 298294 304358 298350
rect 304414 298294 304482 298350
rect 304538 298294 335078 298350
rect 335134 298294 335202 298350
rect 335258 298294 365798 298350
rect 365854 298294 365922 298350
rect 365978 298294 396518 298350
rect 396574 298294 396642 298350
rect 396698 298294 427238 298350
rect 427294 298294 427362 298350
rect 427418 298294 457958 298350
rect 458014 298294 458082 298350
rect 458138 298294 488678 298350
rect 488734 298294 488802 298350
rect 488858 298294 519398 298350
rect 519454 298294 519522 298350
rect 519578 298294 550118 298350
rect 550174 298294 550242 298350
rect 550298 298294 592914 298350
rect 592970 298294 593038 298350
rect 593094 298294 593162 298350
rect 593218 298294 593286 298350
rect 593342 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect -1916 298226 597980 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 27878 298226
rect 27934 298170 28002 298226
rect 28058 298170 58598 298226
rect 58654 298170 58722 298226
rect 58778 298170 89318 298226
rect 89374 298170 89442 298226
rect 89498 298170 120038 298226
rect 120094 298170 120162 298226
rect 120218 298170 150758 298226
rect 150814 298170 150882 298226
rect 150938 298170 181478 298226
rect 181534 298170 181602 298226
rect 181658 298170 212198 298226
rect 212254 298170 212322 298226
rect 212378 298170 242918 298226
rect 242974 298170 243042 298226
rect 243098 298170 273638 298226
rect 273694 298170 273762 298226
rect 273818 298170 304358 298226
rect 304414 298170 304482 298226
rect 304538 298170 335078 298226
rect 335134 298170 335202 298226
rect 335258 298170 365798 298226
rect 365854 298170 365922 298226
rect 365978 298170 396518 298226
rect 396574 298170 396642 298226
rect 396698 298170 427238 298226
rect 427294 298170 427362 298226
rect 427418 298170 457958 298226
rect 458014 298170 458082 298226
rect 458138 298170 488678 298226
rect 488734 298170 488802 298226
rect 488858 298170 519398 298226
rect 519454 298170 519522 298226
rect 519578 298170 550118 298226
rect 550174 298170 550242 298226
rect 550298 298170 592914 298226
rect 592970 298170 593038 298226
rect 593094 298170 593162 298226
rect 593218 298170 593286 298226
rect 593342 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect -1916 298102 597980 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 27878 298102
rect 27934 298046 28002 298102
rect 28058 298046 58598 298102
rect 58654 298046 58722 298102
rect 58778 298046 89318 298102
rect 89374 298046 89442 298102
rect 89498 298046 120038 298102
rect 120094 298046 120162 298102
rect 120218 298046 150758 298102
rect 150814 298046 150882 298102
rect 150938 298046 181478 298102
rect 181534 298046 181602 298102
rect 181658 298046 212198 298102
rect 212254 298046 212322 298102
rect 212378 298046 242918 298102
rect 242974 298046 243042 298102
rect 243098 298046 273638 298102
rect 273694 298046 273762 298102
rect 273818 298046 304358 298102
rect 304414 298046 304482 298102
rect 304538 298046 335078 298102
rect 335134 298046 335202 298102
rect 335258 298046 365798 298102
rect 365854 298046 365922 298102
rect 365978 298046 396518 298102
rect 396574 298046 396642 298102
rect 396698 298046 427238 298102
rect 427294 298046 427362 298102
rect 427418 298046 457958 298102
rect 458014 298046 458082 298102
rect 458138 298046 488678 298102
rect 488734 298046 488802 298102
rect 488858 298046 519398 298102
rect 519454 298046 519522 298102
rect 519578 298046 550118 298102
rect 550174 298046 550242 298102
rect 550298 298046 592914 298102
rect 592970 298046 593038 298102
rect 593094 298046 593162 298102
rect 593218 298046 593286 298102
rect 593342 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect -1916 297978 597980 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 27878 297978
rect 27934 297922 28002 297978
rect 28058 297922 58598 297978
rect 58654 297922 58722 297978
rect 58778 297922 89318 297978
rect 89374 297922 89442 297978
rect 89498 297922 120038 297978
rect 120094 297922 120162 297978
rect 120218 297922 150758 297978
rect 150814 297922 150882 297978
rect 150938 297922 181478 297978
rect 181534 297922 181602 297978
rect 181658 297922 212198 297978
rect 212254 297922 212322 297978
rect 212378 297922 242918 297978
rect 242974 297922 243042 297978
rect 243098 297922 273638 297978
rect 273694 297922 273762 297978
rect 273818 297922 304358 297978
rect 304414 297922 304482 297978
rect 304538 297922 335078 297978
rect 335134 297922 335202 297978
rect 335258 297922 365798 297978
rect 365854 297922 365922 297978
rect 365978 297922 396518 297978
rect 396574 297922 396642 297978
rect 396698 297922 427238 297978
rect 427294 297922 427362 297978
rect 427418 297922 457958 297978
rect 458014 297922 458082 297978
rect 458138 297922 488678 297978
rect 488734 297922 488802 297978
rect 488858 297922 519398 297978
rect 519454 297922 519522 297978
rect 519578 297922 550118 297978
rect 550174 297922 550242 297978
rect 550298 297922 592914 297978
rect 592970 297922 593038 297978
rect 593094 297922 593162 297978
rect 593218 297922 593286 297978
rect 593342 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect -1916 297826 597980 297922
rect -1916 292350 597980 292446
rect -1916 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 5514 292350
rect 5570 292294 5638 292350
rect 5694 292294 5762 292350
rect 5818 292294 5886 292350
rect 5942 292294 12518 292350
rect 12574 292294 12642 292350
rect 12698 292294 43238 292350
rect 43294 292294 43362 292350
rect 43418 292294 73958 292350
rect 74014 292294 74082 292350
rect 74138 292294 104678 292350
rect 104734 292294 104802 292350
rect 104858 292294 135398 292350
rect 135454 292294 135522 292350
rect 135578 292294 166118 292350
rect 166174 292294 166242 292350
rect 166298 292294 196838 292350
rect 196894 292294 196962 292350
rect 197018 292294 227558 292350
rect 227614 292294 227682 292350
rect 227738 292294 258278 292350
rect 258334 292294 258402 292350
rect 258458 292294 288998 292350
rect 289054 292294 289122 292350
rect 289178 292294 319718 292350
rect 319774 292294 319842 292350
rect 319898 292294 350438 292350
rect 350494 292294 350562 292350
rect 350618 292294 381158 292350
rect 381214 292294 381282 292350
rect 381338 292294 411878 292350
rect 411934 292294 412002 292350
rect 412058 292294 442598 292350
rect 442654 292294 442722 292350
rect 442778 292294 473318 292350
rect 473374 292294 473442 292350
rect 473498 292294 504038 292350
rect 504094 292294 504162 292350
rect 504218 292294 534758 292350
rect 534814 292294 534882 292350
rect 534938 292294 565478 292350
rect 565534 292294 565602 292350
rect 565658 292294 589194 292350
rect 589250 292294 589318 292350
rect 589374 292294 589442 292350
rect 589498 292294 589566 292350
rect 589622 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597980 292350
rect -1916 292226 597980 292294
rect -1916 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 5514 292226
rect 5570 292170 5638 292226
rect 5694 292170 5762 292226
rect 5818 292170 5886 292226
rect 5942 292170 12518 292226
rect 12574 292170 12642 292226
rect 12698 292170 43238 292226
rect 43294 292170 43362 292226
rect 43418 292170 73958 292226
rect 74014 292170 74082 292226
rect 74138 292170 104678 292226
rect 104734 292170 104802 292226
rect 104858 292170 135398 292226
rect 135454 292170 135522 292226
rect 135578 292170 166118 292226
rect 166174 292170 166242 292226
rect 166298 292170 196838 292226
rect 196894 292170 196962 292226
rect 197018 292170 227558 292226
rect 227614 292170 227682 292226
rect 227738 292170 258278 292226
rect 258334 292170 258402 292226
rect 258458 292170 288998 292226
rect 289054 292170 289122 292226
rect 289178 292170 319718 292226
rect 319774 292170 319842 292226
rect 319898 292170 350438 292226
rect 350494 292170 350562 292226
rect 350618 292170 381158 292226
rect 381214 292170 381282 292226
rect 381338 292170 411878 292226
rect 411934 292170 412002 292226
rect 412058 292170 442598 292226
rect 442654 292170 442722 292226
rect 442778 292170 473318 292226
rect 473374 292170 473442 292226
rect 473498 292170 504038 292226
rect 504094 292170 504162 292226
rect 504218 292170 534758 292226
rect 534814 292170 534882 292226
rect 534938 292170 565478 292226
rect 565534 292170 565602 292226
rect 565658 292170 589194 292226
rect 589250 292170 589318 292226
rect 589374 292170 589442 292226
rect 589498 292170 589566 292226
rect 589622 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597980 292226
rect -1916 292102 597980 292170
rect -1916 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 5514 292102
rect 5570 292046 5638 292102
rect 5694 292046 5762 292102
rect 5818 292046 5886 292102
rect 5942 292046 12518 292102
rect 12574 292046 12642 292102
rect 12698 292046 43238 292102
rect 43294 292046 43362 292102
rect 43418 292046 73958 292102
rect 74014 292046 74082 292102
rect 74138 292046 104678 292102
rect 104734 292046 104802 292102
rect 104858 292046 135398 292102
rect 135454 292046 135522 292102
rect 135578 292046 166118 292102
rect 166174 292046 166242 292102
rect 166298 292046 196838 292102
rect 196894 292046 196962 292102
rect 197018 292046 227558 292102
rect 227614 292046 227682 292102
rect 227738 292046 258278 292102
rect 258334 292046 258402 292102
rect 258458 292046 288998 292102
rect 289054 292046 289122 292102
rect 289178 292046 319718 292102
rect 319774 292046 319842 292102
rect 319898 292046 350438 292102
rect 350494 292046 350562 292102
rect 350618 292046 381158 292102
rect 381214 292046 381282 292102
rect 381338 292046 411878 292102
rect 411934 292046 412002 292102
rect 412058 292046 442598 292102
rect 442654 292046 442722 292102
rect 442778 292046 473318 292102
rect 473374 292046 473442 292102
rect 473498 292046 504038 292102
rect 504094 292046 504162 292102
rect 504218 292046 534758 292102
rect 534814 292046 534882 292102
rect 534938 292046 565478 292102
rect 565534 292046 565602 292102
rect 565658 292046 589194 292102
rect 589250 292046 589318 292102
rect 589374 292046 589442 292102
rect 589498 292046 589566 292102
rect 589622 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597980 292102
rect -1916 291978 597980 292046
rect -1916 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 5514 291978
rect 5570 291922 5638 291978
rect 5694 291922 5762 291978
rect 5818 291922 5886 291978
rect 5942 291922 12518 291978
rect 12574 291922 12642 291978
rect 12698 291922 43238 291978
rect 43294 291922 43362 291978
rect 43418 291922 73958 291978
rect 74014 291922 74082 291978
rect 74138 291922 104678 291978
rect 104734 291922 104802 291978
rect 104858 291922 135398 291978
rect 135454 291922 135522 291978
rect 135578 291922 166118 291978
rect 166174 291922 166242 291978
rect 166298 291922 196838 291978
rect 196894 291922 196962 291978
rect 197018 291922 227558 291978
rect 227614 291922 227682 291978
rect 227738 291922 258278 291978
rect 258334 291922 258402 291978
rect 258458 291922 288998 291978
rect 289054 291922 289122 291978
rect 289178 291922 319718 291978
rect 319774 291922 319842 291978
rect 319898 291922 350438 291978
rect 350494 291922 350562 291978
rect 350618 291922 381158 291978
rect 381214 291922 381282 291978
rect 381338 291922 411878 291978
rect 411934 291922 412002 291978
rect 412058 291922 442598 291978
rect 442654 291922 442722 291978
rect 442778 291922 473318 291978
rect 473374 291922 473442 291978
rect 473498 291922 504038 291978
rect 504094 291922 504162 291978
rect 504218 291922 534758 291978
rect 534814 291922 534882 291978
rect 534938 291922 565478 291978
rect 565534 291922 565602 291978
rect 565658 291922 589194 291978
rect 589250 291922 589318 291978
rect 589374 291922 589442 291978
rect 589498 291922 589566 291978
rect 589622 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597980 291978
rect -1916 291826 597980 291922
rect -1916 280350 597980 280446
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 27878 280350
rect 27934 280294 28002 280350
rect 28058 280294 58598 280350
rect 58654 280294 58722 280350
rect 58778 280294 89318 280350
rect 89374 280294 89442 280350
rect 89498 280294 120038 280350
rect 120094 280294 120162 280350
rect 120218 280294 150758 280350
rect 150814 280294 150882 280350
rect 150938 280294 181478 280350
rect 181534 280294 181602 280350
rect 181658 280294 212198 280350
rect 212254 280294 212322 280350
rect 212378 280294 242918 280350
rect 242974 280294 243042 280350
rect 243098 280294 273638 280350
rect 273694 280294 273762 280350
rect 273818 280294 304358 280350
rect 304414 280294 304482 280350
rect 304538 280294 335078 280350
rect 335134 280294 335202 280350
rect 335258 280294 365798 280350
rect 365854 280294 365922 280350
rect 365978 280294 396518 280350
rect 396574 280294 396642 280350
rect 396698 280294 427238 280350
rect 427294 280294 427362 280350
rect 427418 280294 457958 280350
rect 458014 280294 458082 280350
rect 458138 280294 488678 280350
rect 488734 280294 488802 280350
rect 488858 280294 519398 280350
rect 519454 280294 519522 280350
rect 519578 280294 550118 280350
rect 550174 280294 550242 280350
rect 550298 280294 592914 280350
rect 592970 280294 593038 280350
rect 593094 280294 593162 280350
rect 593218 280294 593286 280350
rect 593342 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect -1916 280226 597980 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 27878 280226
rect 27934 280170 28002 280226
rect 28058 280170 58598 280226
rect 58654 280170 58722 280226
rect 58778 280170 89318 280226
rect 89374 280170 89442 280226
rect 89498 280170 120038 280226
rect 120094 280170 120162 280226
rect 120218 280170 150758 280226
rect 150814 280170 150882 280226
rect 150938 280170 181478 280226
rect 181534 280170 181602 280226
rect 181658 280170 212198 280226
rect 212254 280170 212322 280226
rect 212378 280170 242918 280226
rect 242974 280170 243042 280226
rect 243098 280170 273638 280226
rect 273694 280170 273762 280226
rect 273818 280170 304358 280226
rect 304414 280170 304482 280226
rect 304538 280170 335078 280226
rect 335134 280170 335202 280226
rect 335258 280170 365798 280226
rect 365854 280170 365922 280226
rect 365978 280170 396518 280226
rect 396574 280170 396642 280226
rect 396698 280170 427238 280226
rect 427294 280170 427362 280226
rect 427418 280170 457958 280226
rect 458014 280170 458082 280226
rect 458138 280170 488678 280226
rect 488734 280170 488802 280226
rect 488858 280170 519398 280226
rect 519454 280170 519522 280226
rect 519578 280170 550118 280226
rect 550174 280170 550242 280226
rect 550298 280170 592914 280226
rect 592970 280170 593038 280226
rect 593094 280170 593162 280226
rect 593218 280170 593286 280226
rect 593342 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect -1916 280102 597980 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 27878 280102
rect 27934 280046 28002 280102
rect 28058 280046 58598 280102
rect 58654 280046 58722 280102
rect 58778 280046 89318 280102
rect 89374 280046 89442 280102
rect 89498 280046 120038 280102
rect 120094 280046 120162 280102
rect 120218 280046 150758 280102
rect 150814 280046 150882 280102
rect 150938 280046 181478 280102
rect 181534 280046 181602 280102
rect 181658 280046 212198 280102
rect 212254 280046 212322 280102
rect 212378 280046 242918 280102
rect 242974 280046 243042 280102
rect 243098 280046 273638 280102
rect 273694 280046 273762 280102
rect 273818 280046 304358 280102
rect 304414 280046 304482 280102
rect 304538 280046 335078 280102
rect 335134 280046 335202 280102
rect 335258 280046 365798 280102
rect 365854 280046 365922 280102
rect 365978 280046 396518 280102
rect 396574 280046 396642 280102
rect 396698 280046 427238 280102
rect 427294 280046 427362 280102
rect 427418 280046 457958 280102
rect 458014 280046 458082 280102
rect 458138 280046 488678 280102
rect 488734 280046 488802 280102
rect 488858 280046 519398 280102
rect 519454 280046 519522 280102
rect 519578 280046 550118 280102
rect 550174 280046 550242 280102
rect 550298 280046 592914 280102
rect 592970 280046 593038 280102
rect 593094 280046 593162 280102
rect 593218 280046 593286 280102
rect 593342 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect -1916 279978 597980 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 27878 279978
rect 27934 279922 28002 279978
rect 28058 279922 58598 279978
rect 58654 279922 58722 279978
rect 58778 279922 89318 279978
rect 89374 279922 89442 279978
rect 89498 279922 120038 279978
rect 120094 279922 120162 279978
rect 120218 279922 150758 279978
rect 150814 279922 150882 279978
rect 150938 279922 181478 279978
rect 181534 279922 181602 279978
rect 181658 279922 212198 279978
rect 212254 279922 212322 279978
rect 212378 279922 242918 279978
rect 242974 279922 243042 279978
rect 243098 279922 273638 279978
rect 273694 279922 273762 279978
rect 273818 279922 304358 279978
rect 304414 279922 304482 279978
rect 304538 279922 335078 279978
rect 335134 279922 335202 279978
rect 335258 279922 365798 279978
rect 365854 279922 365922 279978
rect 365978 279922 396518 279978
rect 396574 279922 396642 279978
rect 396698 279922 427238 279978
rect 427294 279922 427362 279978
rect 427418 279922 457958 279978
rect 458014 279922 458082 279978
rect 458138 279922 488678 279978
rect 488734 279922 488802 279978
rect 488858 279922 519398 279978
rect 519454 279922 519522 279978
rect 519578 279922 550118 279978
rect 550174 279922 550242 279978
rect 550298 279922 592914 279978
rect 592970 279922 593038 279978
rect 593094 279922 593162 279978
rect 593218 279922 593286 279978
rect 593342 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect -1916 279826 597980 279922
rect -1916 274350 597980 274446
rect -1916 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 5514 274350
rect 5570 274294 5638 274350
rect 5694 274294 5762 274350
rect 5818 274294 5886 274350
rect 5942 274294 12518 274350
rect 12574 274294 12642 274350
rect 12698 274294 43238 274350
rect 43294 274294 43362 274350
rect 43418 274294 73958 274350
rect 74014 274294 74082 274350
rect 74138 274294 104678 274350
rect 104734 274294 104802 274350
rect 104858 274294 135398 274350
rect 135454 274294 135522 274350
rect 135578 274294 166118 274350
rect 166174 274294 166242 274350
rect 166298 274294 196838 274350
rect 196894 274294 196962 274350
rect 197018 274294 227558 274350
rect 227614 274294 227682 274350
rect 227738 274294 258278 274350
rect 258334 274294 258402 274350
rect 258458 274294 288998 274350
rect 289054 274294 289122 274350
rect 289178 274294 319718 274350
rect 319774 274294 319842 274350
rect 319898 274294 350438 274350
rect 350494 274294 350562 274350
rect 350618 274294 381158 274350
rect 381214 274294 381282 274350
rect 381338 274294 411878 274350
rect 411934 274294 412002 274350
rect 412058 274294 442598 274350
rect 442654 274294 442722 274350
rect 442778 274294 473318 274350
rect 473374 274294 473442 274350
rect 473498 274294 504038 274350
rect 504094 274294 504162 274350
rect 504218 274294 534758 274350
rect 534814 274294 534882 274350
rect 534938 274294 565478 274350
rect 565534 274294 565602 274350
rect 565658 274294 589194 274350
rect 589250 274294 589318 274350
rect 589374 274294 589442 274350
rect 589498 274294 589566 274350
rect 589622 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597980 274350
rect -1916 274226 597980 274294
rect -1916 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 5514 274226
rect 5570 274170 5638 274226
rect 5694 274170 5762 274226
rect 5818 274170 5886 274226
rect 5942 274170 12518 274226
rect 12574 274170 12642 274226
rect 12698 274170 43238 274226
rect 43294 274170 43362 274226
rect 43418 274170 73958 274226
rect 74014 274170 74082 274226
rect 74138 274170 104678 274226
rect 104734 274170 104802 274226
rect 104858 274170 135398 274226
rect 135454 274170 135522 274226
rect 135578 274170 166118 274226
rect 166174 274170 166242 274226
rect 166298 274170 196838 274226
rect 196894 274170 196962 274226
rect 197018 274170 227558 274226
rect 227614 274170 227682 274226
rect 227738 274170 258278 274226
rect 258334 274170 258402 274226
rect 258458 274170 288998 274226
rect 289054 274170 289122 274226
rect 289178 274170 319718 274226
rect 319774 274170 319842 274226
rect 319898 274170 350438 274226
rect 350494 274170 350562 274226
rect 350618 274170 381158 274226
rect 381214 274170 381282 274226
rect 381338 274170 411878 274226
rect 411934 274170 412002 274226
rect 412058 274170 442598 274226
rect 442654 274170 442722 274226
rect 442778 274170 473318 274226
rect 473374 274170 473442 274226
rect 473498 274170 504038 274226
rect 504094 274170 504162 274226
rect 504218 274170 534758 274226
rect 534814 274170 534882 274226
rect 534938 274170 565478 274226
rect 565534 274170 565602 274226
rect 565658 274170 589194 274226
rect 589250 274170 589318 274226
rect 589374 274170 589442 274226
rect 589498 274170 589566 274226
rect 589622 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597980 274226
rect -1916 274102 597980 274170
rect -1916 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 5514 274102
rect 5570 274046 5638 274102
rect 5694 274046 5762 274102
rect 5818 274046 5886 274102
rect 5942 274046 12518 274102
rect 12574 274046 12642 274102
rect 12698 274046 43238 274102
rect 43294 274046 43362 274102
rect 43418 274046 73958 274102
rect 74014 274046 74082 274102
rect 74138 274046 104678 274102
rect 104734 274046 104802 274102
rect 104858 274046 135398 274102
rect 135454 274046 135522 274102
rect 135578 274046 166118 274102
rect 166174 274046 166242 274102
rect 166298 274046 196838 274102
rect 196894 274046 196962 274102
rect 197018 274046 227558 274102
rect 227614 274046 227682 274102
rect 227738 274046 258278 274102
rect 258334 274046 258402 274102
rect 258458 274046 288998 274102
rect 289054 274046 289122 274102
rect 289178 274046 319718 274102
rect 319774 274046 319842 274102
rect 319898 274046 350438 274102
rect 350494 274046 350562 274102
rect 350618 274046 381158 274102
rect 381214 274046 381282 274102
rect 381338 274046 411878 274102
rect 411934 274046 412002 274102
rect 412058 274046 442598 274102
rect 442654 274046 442722 274102
rect 442778 274046 473318 274102
rect 473374 274046 473442 274102
rect 473498 274046 504038 274102
rect 504094 274046 504162 274102
rect 504218 274046 534758 274102
rect 534814 274046 534882 274102
rect 534938 274046 565478 274102
rect 565534 274046 565602 274102
rect 565658 274046 589194 274102
rect 589250 274046 589318 274102
rect 589374 274046 589442 274102
rect 589498 274046 589566 274102
rect 589622 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597980 274102
rect -1916 273978 597980 274046
rect -1916 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 5514 273978
rect 5570 273922 5638 273978
rect 5694 273922 5762 273978
rect 5818 273922 5886 273978
rect 5942 273922 12518 273978
rect 12574 273922 12642 273978
rect 12698 273922 43238 273978
rect 43294 273922 43362 273978
rect 43418 273922 73958 273978
rect 74014 273922 74082 273978
rect 74138 273922 104678 273978
rect 104734 273922 104802 273978
rect 104858 273922 135398 273978
rect 135454 273922 135522 273978
rect 135578 273922 166118 273978
rect 166174 273922 166242 273978
rect 166298 273922 196838 273978
rect 196894 273922 196962 273978
rect 197018 273922 227558 273978
rect 227614 273922 227682 273978
rect 227738 273922 258278 273978
rect 258334 273922 258402 273978
rect 258458 273922 288998 273978
rect 289054 273922 289122 273978
rect 289178 273922 319718 273978
rect 319774 273922 319842 273978
rect 319898 273922 350438 273978
rect 350494 273922 350562 273978
rect 350618 273922 381158 273978
rect 381214 273922 381282 273978
rect 381338 273922 411878 273978
rect 411934 273922 412002 273978
rect 412058 273922 442598 273978
rect 442654 273922 442722 273978
rect 442778 273922 473318 273978
rect 473374 273922 473442 273978
rect 473498 273922 504038 273978
rect 504094 273922 504162 273978
rect 504218 273922 534758 273978
rect 534814 273922 534882 273978
rect 534938 273922 565478 273978
rect 565534 273922 565602 273978
rect 565658 273922 589194 273978
rect 589250 273922 589318 273978
rect 589374 273922 589442 273978
rect 589498 273922 589566 273978
rect 589622 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597980 273978
rect -1916 273826 597980 273922
rect -1916 262350 597980 262446
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 27878 262350
rect 27934 262294 28002 262350
rect 28058 262294 58598 262350
rect 58654 262294 58722 262350
rect 58778 262294 89318 262350
rect 89374 262294 89442 262350
rect 89498 262294 120038 262350
rect 120094 262294 120162 262350
rect 120218 262294 150758 262350
rect 150814 262294 150882 262350
rect 150938 262294 181478 262350
rect 181534 262294 181602 262350
rect 181658 262294 212198 262350
rect 212254 262294 212322 262350
rect 212378 262294 242918 262350
rect 242974 262294 243042 262350
rect 243098 262294 273638 262350
rect 273694 262294 273762 262350
rect 273818 262294 304358 262350
rect 304414 262294 304482 262350
rect 304538 262294 335078 262350
rect 335134 262294 335202 262350
rect 335258 262294 365798 262350
rect 365854 262294 365922 262350
rect 365978 262294 396518 262350
rect 396574 262294 396642 262350
rect 396698 262294 427238 262350
rect 427294 262294 427362 262350
rect 427418 262294 457958 262350
rect 458014 262294 458082 262350
rect 458138 262294 488678 262350
rect 488734 262294 488802 262350
rect 488858 262294 519398 262350
rect 519454 262294 519522 262350
rect 519578 262294 550118 262350
rect 550174 262294 550242 262350
rect 550298 262294 592914 262350
rect 592970 262294 593038 262350
rect 593094 262294 593162 262350
rect 593218 262294 593286 262350
rect 593342 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect -1916 262226 597980 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 27878 262226
rect 27934 262170 28002 262226
rect 28058 262170 58598 262226
rect 58654 262170 58722 262226
rect 58778 262170 89318 262226
rect 89374 262170 89442 262226
rect 89498 262170 120038 262226
rect 120094 262170 120162 262226
rect 120218 262170 150758 262226
rect 150814 262170 150882 262226
rect 150938 262170 181478 262226
rect 181534 262170 181602 262226
rect 181658 262170 212198 262226
rect 212254 262170 212322 262226
rect 212378 262170 242918 262226
rect 242974 262170 243042 262226
rect 243098 262170 273638 262226
rect 273694 262170 273762 262226
rect 273818 262170 304358 262226
rect 304414 262170 304482 262226
rect 304538 262170 335078 262226
rect 335134 262170 335202 262226
rect 335258 262170 365798 262226
rect 365854 262170 365922 262226
rect 365978 262170 396518 262226
rect 396574 262170 396642 262226
rect 396698 262170 427238 262226
rect 427294 262170 427362 262226
rect 427418 262170 457958 262226
rect 458014 262170 458082 262226
rect 458138 262170 488678 262226
rect 488734 262170 488802 262226
rect 488858 262170 519398 262226
rect 519454 262170 519522 262226
rect 519578 262170 550118 262226
rect 550174 262170 550242 262226
rect 550298 262170 592914 262226
rect 592970 262170 593038 262226
rect 593094 262170 593162 262226
rect 593218 262170 593286 262226
rect 593342 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect -1916 262102 597980 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 27878 262102
rect 27934 262046 28002 262102
rect 28058 262046 58598 262102
rect 58654 262046 58722 262102
rect 58778 262046 89318 262102
rect 89374 262046 89442 262102
rect 89498 262046 120038 262102
rect 120094 262046 120162 262102
rect 120218 262046 150758 262102
rect 150814 262046 150882 262102
rect 150938 262046 181478 262102
rect 181534 262046 181602 262102
rect 181658 262046 212198 262102
rect 212254 262046 212322 262102
rect 212378 262046 242918 262102
rect 242974 262046 243042 262102
rect 243098 262046 273638 262102
rect 273694 262046 273762 262102
rect 273818 262046 304358 262102
rect 304414 262046 304482 262102
rect 304538 262046 335078 262102
rect 335134 262046 335202 262102
rect 335258 262046 365798 262102
rect 365854 262046 365922 262102
rect 365978 262046 396518 262102
rect 396574 262046 396642 262102
rect 396698 262046 427238 262102
rect 427294 262046 427362 262102
rect 427418 262046 457958 262102
rect 458014 262046 458082 262102
rect 458138 262046 488678 262102
rect 488734 262046 488802 262102
rect 488858 262046 519398 262102
rect 519454 262046 519522 262102
rect 519578 262046 550118 262102
rect 550174 262046 550242 262102
rect 550298 262046 592914 262102
rect 592970 262046 593038 262102
rect 593094 262046 593162 262102
rect 593218 262046 593286 262102
rect 593342 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect -1916 261978 597980 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 27878 261978
rect 27934 261922 28002 261978
rect 28058 261922 58598 261978
rect 58654 261922 58722 261978
rect 58778 261922 89318 261978
rect 89374 261922 89442 261978
rect 89498 261922 120038 261978
rect 120094 261922 120162 261978
rect 120218 261922 150758 261978
rect 150814 261922 150882 261978
rect 150938 261922 181478 261978
rect 181534 261922 181602 261978
rect 181658 261922 212198 261978
rect 212254 261922 212322 261978
rect 212378 261922 242918 261978
rect 242974 261922 243042 261978
rect 243098 261922 273638 261978
rect 273694 261922 273762 261978
rect 273818 261922 304358 261978
rect 304414 261922 304482 261978
rect 304538 261922 335078 261978
rect 335134 261922 335202 261978
rect 335258 261922 365798 261978
rect 365854 261922 365922 261978
rect 365978 261922 396518 261978
rect 396574 261922 396642 261978
rect 396698 261922 427238 261978
rect 427294 261922 427362 261978
rect 427418 261922 457958 261978
rect 458014 261922 458082 261978
rect 458138 261922 488678 261978
rect 488734 261922 488802 261978
rect 488858 261922 519398 261978
rect 519454 261922 519522 261978
rect 519578 261922 550118 261978
rect 550174 261922 550242 261978
rect 550298 261922 592914 261978
rect 592970 261922 593038 261978
rect 593094 261922 593162 261978
rect 593218 261922 593286 261978
rect 593342 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect -1916 261826 597980 261922
rect -1916 256350 597980 256446
rect -1916 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 5514 256350
rect 5570 256294 5638 256350
rect 5694 256294 5762 256350
rect 5818 256294 5886 256350
rect 5942 256294 12518 256350
rect 12574 256294 12642 256350
rect 12698 256294 43238 256350
rect 43294 256294 43362 256350
rect 43418 256294 73958 256350
rect 74014 256294 74082 256350
rect 74138 256294 104678 256350
rect 104734 256294 104802 256350
rect 104858 256294 135398 256350
rect 135454 256294 135522 256350
rect 135578 256294 166118 256350
rect 166174 256294 166242 256350
rect 166298 256294 196838 256350
rect 196894 256294 196962 256350
rect 197018 256294 227558 256350
rect 227614 256294 227682 256350
rect 227738 256294 258278 256350
rect 258334 256294 258402 256350
rect 258458 256294 288998 256350
rect 289054 256294 289122 256350
rect 289178 256294 319718 256350
rect 319774 256294 319842 256350
rect 319898 256294 350438 256350
rect 350494 256294 350562 256350
rect 350618 256294 381158 256350
rect 381214 256294 381282 256350
rect 381338 256294 411878 256350
rect 411934 256294 412002 256350
rect 412058 256294 442598 256350
rect 442654 256294 442722 256350
rect 442778 256294 473318 256350
rect 473374 256294 473442 256350
rect 473498 256294 504038 256350
rect 504094 256294 504162 256350
rect 504218 256294 534758 256350
rect 534814 256294 534882 256350
rect 534938 256294 565478 256350
rect 565534 256294 565602 256350
rect 565658 256294 589194 256350
rect 589250 256294 589318 256350
rect 589374 256294 589442 256350
rect 589498 256294 589566 256350
rect 589622 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597980 256350
rect -1916 256226 597980 256294
rect -1916 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 5514 256226
rect 5570 256170 5638 256226
rect 5694 256170 5762 256226
rect 5818 256170 5886 256226
rect 5942 256170 12518 256226
rect 12574 256170 12642 256226
rect 12698 256170 43238 256226
rect 43294 256170 43362 256226
rect 43418 256170 73958 256226
rect 74014 256170 74082 256226
rect 74138 256170 104678 256226
rect 104734 256170 104802 256226
rect 104858 256170 135398 256226
rect 135454 256170 135522 256226
rect 135578 256170 166118 256226
rect 166174 256170 166242 256226
rect 166298 256170 196838 256226
rect 196894 256170 196962 256226
rect 197018 256170 227558 256226
rect 227614 256170 227682 256226
rect 227738 256170 258278 256226
rect 258334 256170 258402 256226
rect 258458 256170 288998 256226
rect 289054 256170 289122 256226
rect 289178 256170 319718 256226
rect 319774 256170 319842 256226
rect 319898 256170 350438 256226
rect 350494 256170 350562 256226
rect 350618 256170 381158 256226
rect 381214 256170 381282 256226
rect 381338 256170 411878 256226
rect 411934 256170 412002 256226
rect 412058 256170 442598 256226
rect 442654 256170 442722 256226
rect 442778 256170 473318 256226
rect 473374 256170 473442 256226
rect 473498 256170 504038 256226
rect 504094 256170 504162 256226
rect 504218 256170 534758 256226
rect 534814 256170 534882 256226
rect 534938 256170 565478 256226
rect 565534 256170 565602 256226
rect 565658 256170 589194 256226
rect 589250 256170 589318 256226
rect 589374 256170 589442 256226
rect 589498 256170 589566 256226
rect 589622 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597980 256226
rect -1916 256102 597980 256170
rect -1916 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 5514 256102
rect 5570 256046 5638 256102
rect 5694 256046 5762 256102
rect 5818 256046 5886 256102
rect 5942 256046 12518 256102
rect 12574 256046 12642 256102
rect 12698 256046 43238 256102
rect 43294 256046 43362 256102
rect 43418 256046 73958 256102
rect 74014 256046 74082 256102
rect 74138 256046 104678 256102
rect 104734 256046 104802 256102
rect 104858 256046 135398 256102
rect 135454 256046 135522 256102
rect 135578 256046 166118 256102
rect 166174 256046 166242 256102
rect 166298 256046 196838 256102
rect 196894 256046 196962 256102
rect 197018 256046 227558 256102
rect 227614 256046 227682 256102
rect 227738 256046 258278 256102
rect 258334 256046 258402 256102
rect 258458 256046 288998 256102
rect 289054 256046 289122 256102
rect 289178 256046 319718 256102
rect 319774 256046 319842 256102
rect 319898 256046 350438 256102
rect 350494 256046 350562 256102
rect 350618 256046 381158 256102
rect 381214 256046 381282 256102
rect 381338 256046 411878 256102
rect 411934 256046 412002 256102
rect 412058 256046 442598 256102
rect 442654 256046 442722 256102
rect 442778 256046 473318 256102
rect 473374 256046 473442 256102
rect 473498 256046 504038 256102
rect 504094 256046 504162 256102
rect 504218 256046 534758 256102
rect 534814 256046 534882 256102
rect 534938 256046 565478 256102
rect 565534 256046 565602 256102
rect 565658 256046 589194 256102
rect 589250 256046 589318 256102
rect 589374 256046 589442 256102
rect 589498 256046 589566 256102
rect 589622 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597980 256102
rect -1916 255978 597980 256046
rect -1916 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 5514 255978
rect 5570 255922 5638 255978
rect 5694 255922 5762 255978
rect 5818 255922 5886 255978
rect 5942 255922 12518 255978
rect 12574 255922 12642 255978
rect 12698 255922 43238 255978
rect 43294 255922 43362 255978
rect 43418 255922 73958 255978
rect 74014 255922 74082 255978
rect 74138 255922 104678 255978
rect 104734 255922 104802 255978
rect 104858 255922 135398 255978
rect 135454 255922 135522 255978
rect 135578 255922 166118 255978
rect 166174 255922 166242 255978
rect 166298 255922 196838 255978
rect 196894 255922 196962 255978
rect 197018 255922 227558 255978
rect 227614 255922 227682 255978
rect 227738 255922 258278 255978
rect 258334 255922 258402 255978
rect 258458 255922 288998 255978
rect 289054 255922 289122 255978
rect 289178 255922 319718 255978
rect 319774 255922 319842 255978
rect 319898 255922 350438 255978
rect 350494 255922 350562 255978
rect 350618 255922 381158 255978
rect 381214 255922 381282 255978
rect 381338 255922 411878 255978
rect 411934 255922 412002 255978
rect 412058 255922 442598 255978
rect 442654 255922 442722 255978
rect 442778 255922 473318 255978
rect 473374 255922 473442 255978
rect 473498 255922 504038 255978
rect 504094 255922 504162 255978
rect 504218 255922 534758 255978
rect 534814 255922 534882 255978
rect 534938 255922 565478 255978
rect 565534 255922 565602 255978
rect 565658 255922 589194 255978
rect 589250 255922 589318 255978
rect 589374 255922 589442 255978
rect 589498 255922 589566 255978
rect 589622 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597980 255978
rect -1916 255826 597980 255922
rect -1916 244350 597980 244446
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 27878 244350
rect 27934 244294 28002 244350
rect 28058 244294 58598 244350
rect 58654 244294 58722 244350
rect 58778 244294 89318 244350
rect 89374 244294 89442 244350
rect 89498 244294 120038 244350
rect 120094 244294 120162 244350
rect 120218 244294 150758 244350
rect 150814 244294 150882 244350
rect 150938 244294 181478 244350
rect 181534 244294 181602 244350
rect 181658 244294 212198 244350
rect 212254 244294 212322 244350
rect 212378 244294 242918 244350
rect 242974 244294 243042 244350
rect 243098 244294 273638 244350
rect 273694 244294 273762 244350
rect 273818 244294 304358 244350
rect 304414 244294 304482 244350
rect 304538 244294 335078 244350
rect 335134 244294 335202 244350
rect 335258 244294 365798 244350
rect 365854 244294 365922 244350
rect 365978 244294 396518 244350
rect 396574 244294 396642 244350
rect 396698 244294 427238 244350
rect 427294 244294 427362 244350
rect 427418 244294 457958 244350
rect 458014 244294 458082 244350
rect 458138 244294 488678 244350
rect 488734 244294 488802 244350
rect 488858 244294 519398 244350
rect 519454 244294 519522 244350
rect 519578 244294 550118 244350
rect 550174 244294 550242 244350
rect 550298 244294 592914 244350
rect 592970 244294 593038 244350
rect 593094 244294 593162 244350
rect 593218 244294 593286 244350
rect 593342 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect -1916 244226 597980 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 27878 244226
rect 27934 244170 28002 244226
rect 28058 244170 58598 244226
rect 58654 244170 58722 244226
rect 58778 244170 89318 244226
rect 89374 244170 89442 244226
rect 89498 244170 120038 244226
rect 120094 244170 120162 244226
rect 120218 244170 150758 244226
rect 150814 244170 150882 244226
rect 150938 244170 181478 244226
rect 181534 244170 181602 244226
rect 181658 244170 212198 244226
rect 212254 244170 212322 244226
rect 212378 244170 242918 244226
rect 242974 244170 243042 244226
rect 243098 244170 273638 244226
rect 273694 244170 273762 244226
rect 273818 244170 304358 244226
rect 304414 244170 304482 244226
rect 304538 244170 335078 244226
rect 335134 244170 335202 244226
rect 335258 244170 365798 244226
rect 365854 244170 365922 244226
rect 365978 244170 396518 244226
rect 396574 244170 396642 244226
rect 396698 244170 427238 244226
rect 427294 244170 427362 244226
rect 427418 244170 457958 244226
rect 458014 244170 458082 244226
rect 458138 244170 488678 244226
rect 488734 244170 488802 244226
rect 488858 244170 519398 244226
rect 519454 244170 519522 244226
rect 519578 244170 550118 244226
rect 550174 244170 550242 244226
rect 550298 244170 592914 244226
rect 592970 244170 593038 244226
rect 593094 244170 593162 244226
rect 593218 244170 593286 244226
rect 593342 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect -1916 244102 597980 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 27878 244102
rect 27934 244046 28002 244102
rect 28058 244046 58598 244102
rect 58654 244046 58722 244102
rect 58778 244046 89318 244102
rect 89374 244046 89442 244102
rect 89498 244046 120038 244102
rect 120094 244046 120162 244102
rect 120218 244046 150758 244102
rect 150814 244046 150882 244102
rect 150938 244046 181478 244102
rect 181534 244046 181602 244102
rect 181658 244046 212198 244102
rect 212254 244046 212322 244102
rect 212378 244046 242918 244102
rect 242974 244046 243042 244102
rect 243098 244046 273638 244102
rect 273694 244046 273762 244102
rect 273818 244046 304358 244102
rect 304414 244046 304482 244102
rect 304538 244046 335078 244102
rect 335134 244046 335202 244102
rect 335258 244046 365798 244102
rect 365854 244046 365922 244102
rect 365978 244046 396518 244102
rect 396574 244046 396642 244102
rect 396698 244046 427238 244102
rect 427294 244046 427362 244102
rect 427418 244046 457958 244102
rect 458014 244046 458082 244102
rect 458138 244046 488678 244102
rect 488734 244046 488802 244102
rect 488858 244046 519398 244102
rect 519454 244046 519522 244102
rect 519578 244046 550118 244102
rect 550174 244046 550242 244102
rect 550298 244046 592914 244102
rect 592970 244046 593038 244102
rect 593094 244046 593162 244102
rect 593218 244046 593286 244102
rect 593342 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect -1916 243978 597980 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 27878 243978
rect 27934 243922 28002 243978
rect 28058 243922 58598 243978
rect 58654 243922 58722 243978
rect 58778 243922 89318 243978
rect 89374 243922 89442 243978
rect 89498 243922 120038 243978
rect 120094 243922 120162 243978
rect 120218 243922 150758 243978
rect 150814 243922 150882 243978
rect 150938 243922 181478 243978
rect 181534 243922 181602 243978
rect 181658 243922 212198 243978
rect 212254 243922 212322 243978
rect 212378 243922 242918 243978
rect 242974 243922 243042 243978
rect 243098 243922 273638 243978
rect 273694 243922 273762 243978
rect 273818 243922 304358 243978
rect 304414 243922 304482 243978
rect 304538 243922 335078 243978
rect 335134 243922 335202 243978
rect 335258 243922 365798 243978
rect 365854 243922 365922 243978
rect 365978 243922 396518 243978
rect 396574 243922 396642 243978
rect 396698 243922 427238 243978
rect 427294 243922 427362 243978
rect 427418 243922 457958 243978
rect 458014 243922 458082 243978
rect 458138 243922 488678 243978
rect 488734 243922 488802 243978
rect 488858 243922 519398 243978
rect 519454 243922 519522 243978
rect 519578 243922 550118 243978
rect 550174 243922 550242 243978
rect 550298 243922 592914 243978
rect 592970 243922 593038 243978
rect 593094 243922 593162 243978
rect 593218 243922 593286 243978
rect 593342 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect -1916 243826 597980 243922
rect -1916 238350 597980 238446
rect -1916 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 5514 238350
rect 5570 238294 5638 238350
rect 5694 238294 5762 238350
rect 5818 238294 5886 238350
rect 5942 238294 12518 238350
rect 12574 238294 12642 238350
rect 12698 238294 43238 238350
rect 43294 238294 43362 238350
rect 43418 238294 73958 238350
rect 74014 238294 74082 238350
rect 74138 238294 104678 238350
rect 104734 238294 104802 238350
rect 104858 238294 135398 238350
rect 135454 238294 135522 238350
rect 135578 238294 166118 238350
rect 166174 238294 166242 238350
rect 166298 238294 196838 238350
rect 196894 238294 196962 238350
rect 197018 238294 227558 238350
rect 227614 238294 227682 238350
rect 227738 238294 258278 238350
rect 258334 238294 258402 238350
rect 258458 238294 288998 238350
rect 289054 238294 289122 238350
rect 289178 238294 319718 238350
rect 319774 238294 319842 238350
rect 319898 238294 350438 238350
rect 350494 238294 350562 238350
rect 350618 238294 381158 238350
rect 381214 238294 381282 238350
rect 381338 238294 411878 238350
rect 411934 238294 412002 238350
rect 412058 238294 442598 238350
rect 442654 238294 442722 238350
rect 442778 238294 473318 238350
rect 473374 238294 473442 238350
rect 473498 238294 504038 238350
rect 504094 238294 504162 238350
rect 504218 238294 534758 238350
rect 534814 238294 534882 238350
rect 534938 238294 565478 238350
rect 565534 238294 565602 238350
rect 565658 238294 589194 238350
rect 589250 238294 589318 238350
rect 589374 238294 589442 238350
rect 589498 238294 589566 238350
rect 589622 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597980 238350
rect -1916 238226 597980 238294
rect -1916 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 5514 238226
rect 5570 238170 5638 238226
rect 5694 238170 5762 238226
rect 5818 238170 5886 238226
rect 5942 238170 12518 238226
rect 12574 238170 12642 238226
rect 12698 238170 43238 238226
rect 43294 238170 43362 238226
rect 43418 238170 73958 238226
rect 74014 238170 74082 238226
rect 74138 238170 104678 238226
rect 104734 238170 104802 238226
rect 104858 238170 135398 238226
rect 135454 238170 135522 238226
rect 135578 238170 166118 238226
rect 166174 238170 166242 238226
rect 166298 238170 196838 238226
rect 196894 238170 196962 238226
rect 197018 238170 227558 238226
rect 227614 238170 227682 238226
rect 227738 238170 258278 238226
rect 258334 238170 258402 238226
rect 258458 238170 288998 238226
rect 289054 238170 289122 238226
rect 289178 238170 319718 238226
rect 319774 238170 319842 238226
rect 319898 238170 350438 238226
rect 350494 238170 350562 238226
rect 350618 238170 381158 238226
rect 381214 238170 381282 238226
rect 381338 238170 411878 238226
rect 411934 238170 412002 238226
rect 412058 238170 442598 238226
rect 442654 238170 442722 238226
rect 442778 238170 473318 238226
rect 473374 238170 473442 238226
rect 473498 238170 504038 238226
rect 504094 238170 504162 238226
rect 504218 238170 534758 238226
rect 534814 238170 534882 238226
rect 534938 238170 565478 238226
rect 565534 238170 565602 238226
rect 565658 238170 589194 238226
rect 589250 238170 589318 238226
rect 589374 238170 589442 238226
rect 589498 238170 589566 238226
rect 589622 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597980 238226
rect -1916 238102 597980 238170
rect -1916 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 5514 238102
rect 5570 238046 5638 238102
rect 5694 238046 5762 238102
rect 5818 238046 5886 238102
rect 5942 238046 12518 238102
rect 12574 238046 12642 238102
rect 12698 238046 43238 238102
rect 43294 238046 43362 238102
rect 43418 238046 73958 238102
rect 74014 238046 74082 238102
rect 74138 238046 104678 238102
rect 104734 238046 104802 238102
rect 104858 238046 135398 238102
rect 135454 238046 135522 238102
rect 135578 238046 166118 238102
rect 166174 238046 166242 238102
rect 166298 238046 196838 238102
rect 196894 238046 196962 238102
rect 197018 238046 227558 238102
rect 227614 238046 227682 238102
rect 227738 238046 258278 238102
rect 258334 238046 258402 238102
rect 258458 238046 288998 238102
rect 289054 238046 289122 238102
rect 289178 238046 319718 238102
rect 319774 238046 319842 238102
rect 319898 238046 350438 238102
rect 350494 238046 350562 238102
rect 350618 238046 381158 238102
rect 381214 238046 381282 238102
rect 381338 238046 411878 238102
rect 411934 238046 412002 238102
rect 412058 238046 442598 238102
rect 442654 238046 442722 238102
rect 442778 238046 473318 238102
rect 473374 238046 473442 238102
rect 473498 238046 504038 238102
rect 504094 238046 504162 238102
rect 504218 238046 534758 238102
rect 534814 238046 534882 238102
rect 534938 238046 565478 238102
rect 565534 238046 565602 238102
rect 565658 238046 589194 238102
rect 589250 238046 589318 238102
rect 589374 238046 589442 238102
rect 589498 238046 589566 238102
rect 589622 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597980 238102
rect -1916 237978 597980 238046
rect -1916 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 5514 237978
rect 5570 237922 5638 237978
rect 5694 237922 5762 237978
rect 5818 237922 5886 237978
rect 5942 237922 12518 237978
rect 12574 237922 12642 237978
rect 12698 237922 43238 237978
rect 43294 237922 43362 237978
rect 43418 237922 73958 237978
rect 74014 237922 74082 237978
rect 74138 237922 104678 237978
rect 104734 237922 104802 237978
rect 104858 237922 135398 237978
rect 135454 237922 135522 237978
rect 135578 237922 166118 237978
rect 166174 237922 166242 237978
rect 166298 237922 196838 237978
rect 196894 237922 196962 237978
rect 197018 237922 227558 237978
rect 227614 237922 227682 237978
rect 227738 237922 258278 237978
rect 258334 237922 258402 237978
rect 258458 237922 288998 237978
rect 289054 237922 289122 237978
rect 289178 237922 319718 237978
rect 319774 237922 319842 237978
rect 319898 237922 350438 237978
rect 350494 237922 350562 237978
rect 350618 237922 381158 237978
rect 381214 237922 381282 237978
rect 381338 237922 411878 237978
rect 411934 237922 412002 237978
rect 412058 237922 442598 237978
rect 442654 237922 442722 237978
rect 442778 237922 473318 237978
rect 473374 237922 473442 237978
rect 473498 237922 504038 237978
rect 504094 237922 504162 237978
rect 504218 237922 534758 237978
rect 534814 237922 534882 237978
rect 534938 237922 565478 237978
rect 565534 237922 565602 237978
rect 565658 237922 589194 237978
rect 589250 237922 589318 237978
rect 589374 237922 589442 237978
rect 589498 237922 589566 237978
rect 589622 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597980 237978
rect -1916 237826 597980 237922
rect -1916 226350 597980 226446
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 27878 226350
rect 27934 226294 28002 226350
rect 28058 226294 58598 226350
rect 58654 226294 58722 226350
rect 58778 226294 89318 226350
rect 89374 226294 89442 226350
rect 89498 226294 120038 226350
rect 120094 226294 120162 226350
rect 120218 226294 150758 226350
rect 150814 226294 150882 226350
rect 150938 226294 181478 226350
rect 181534 226294 181602 226350
rect 181658 226294 212198 226350
rect 212254 226294 212322 226350
rect 212378 226294 242918 226350
rect 242974 226294 243042 226350
rect 243098 226294 273638 226350
rect 273694 226294 273762 226350
rect 273818 226294 304358 226350
rect 304414 226294 304482 226350
rect 304538 226294 335078 226350
rect 335134 226294 335202 226350
rect 335258 226294 365798 226350
rect 365854 226294 365922 226350
rect 365978 226294 396518 226350
rect 396574 226294 396642 226350
rect 396698 226294 427238 226350
rect 427294 226294 427362 226350
rect 427418 226294 457958 226350
rect 458014 226294 458082 226350
rect 458138 226294 488678 226350
rect 488734 226294 488802 226350
rect 488858 226294 519398 226350
rect 519454 226294 519522 226350
rect 519578 226294 550118 226350
rect 550174 226294 550242 226350
rect 550298 226294 592914 226350
rect 592970 226294 593038 226350
rect 593094 226294 593162 226350
rect 593218 226294 593286 226350
rect 593342 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect -1916 226226 597980 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 27878 226226
rect 27934 226170 28002 226226
rect 28058 226170 58598 226226
rect 58654 226170 58722 226226
rect 58778 226170 89318 226226
rect 89374 226170 89442 226226
rect 89498 226170 120038 226226
rect 120094 226170 120162 226226
rect 120218 226170 150758 226226
rect 150814 226170 150882 226226
rect 150938 226170 181478 226226
rect 181534 226170 181602 226226
rect 181658 226170 212198 226226
rect 212254 226170 212322 226226
rect 212378 226170 242918 226226
rect 242974 226170 243042 226226
rect 243098 226170 273638 226226
rect 273694 226170 273762 226226
rect 273818 226170 304358 226226
rect 304414 226170 304482 226226
rect 304538 226170 335078 226226
rect 335134 226170 335202 226226
rect 335258 226170 365798 226226
rect 365854 226170 365922 226226
rect 365978 226170 396518 226226
rect 396574 226170 396642 226226
rect 396698 226170 427238 226226
rect 427294 226170 427362 226226
rect 427418 226170 457958 226226
rect 458014 226170 458082 226226
rect 458138 226170 488678 226226
rect 488734 226170 488802 226226
rect 488858 226170 519398 226226
rect 519454 226170 519522 226226
rect 519578 226170 550118 226226
rect 550174 226170 550242 226226
rect 550298 226170 592914 226226
rect 592970 226170 593038 226226
rect 593094 226170 593162 226226
rect 593218 226170 593286 226226
rect 593342 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect -1916 226102 597980 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 27878 226102
rect 27934 226046 28002 226102
rect 28058 226046 58598 226102
rect 58654 226046 58722 226102
rect 58778 226046 89318 226102
rect 89374 226046 89442 226102
rect 89498 226046 120038 226102
rect 120094 226046 120162 226102
rect 120218 226046 150758 226102
rect 150814 226046 150882 226102
rect 150938 226046 181478 226102
rect 181534 226046 181602 226102
rect 181658 226046 212198 226102
rect 212254 226046 212322 226102
rect 212378 226046 242918 226102
rect 242974 226046 243042 226102
rect 243098 226046 273638 226102
rect 273694 226046 273762 226102
rect 273818 226046 304358 226102
rect 304414 226046 304482 226102
rect 304538 226046 335078 226102
rect 335134 226046 335202 226102
rect 335258 226046 365798 226102
rect 365854 226046 365922 226102
rect 365978 226046 396518 226102
rect 396574 226046 396642 226102
rect 396698 226046 427238 226102
rect 427294 226046 427362 226102
rect 427418 226046 457958 226102
rect 458014 226046 458082 226102
rect 458138 226046 488678 226102
rect 488734 226046 488802 226102
rect 488858 226046 519398 226102
rect 519454 226046 519522 226102
rect 519578 226046 550118 226102
rect 550174 226046 550242 226102
rect 550298 226046 592914 226102
rect 592970 226046 593038 226102
rect 593094 226046 593162 226102
rect 593218 226046 593286 226102
rect 593342 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect -1916 225978 597980 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 27878 225978
rect 27934 225922 28002 225978
rect 28058 225922 58598 225978
rect 58654 225922 58722 225978
rect 58778 225922 89318 225978
rect 89374 225922 89442 225978
rect 89498 225922 120038 225978
rect 120094 225922 120162 225978
rect 120218 225922 150758 225978
rect 150814 225922 150882 225978
rect 150938 225922 181478 225978
rect 181534 225922 181602 225978
rect 181658 225922 212198 225978
rect 212254 225922 212322 225978
rect 212378 225922 242918 225978
rect 242974 225922 243042 225978
rect 243098 225922 273638 225978
rect 273694 225922 273762 225978
rect 273818 225922 304358 225978
rect 304414 225922 304482 225978
rect 304538 225922 335078 225978
rect 335134 225922 335202 225978
rect 335258 225922 365798 225978
rect 365854 225922 365922 225978
rect 365978 225922 396518 225978
rect 396574 225922 396642 225978
rect 396698 225922 427238 225978
rect 427294 225922 427362 225978
rect 427418 225922 457958 225978
rect 458014 225922 458082 225978
rect 458138 225922 488678 225978
rect 488734 225922 488802 225978
rect 488858 225922 519398 225978
rect 519454 225922 519522 225978
rect 519578 225922 550118 225978
rect 550174 225922 550242 225978
rect 550298 225922 592914 225978
rect 592970 225922 593038 225978
rect 593094 225922 593162 225978
rect 593218 225922 593286 225978
rect 593342 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect -1916 225826 597980 225922
rect -1916 220350 597980 220446
rect -1916 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 5514 220350
rect 5570 220294 5638 220350
rect 5694 220294 5762 220350
rect 5818 220294 5886 220350
rect 5942 220294 12518 220350
rect 12574 220294 12642 220350
rect 12698 220294 43238 220350
rect 43294 220294 43362 220350
rect 43418 220294 73958 220350
rect 74014 220294 74082 220350
rect 74138 220294 104678 220350
rect 104734 220294 104802 220350
rect 104858 220294 135398 220350
rect 135454 220294 135522 220350
rect 135578 220294 166118 220350
rect 166174 220294 166242 220350
rect 166298 220294 196838 220350
rect 196894 220294 196962 220350
rect 197018 220294 227558 220350
rect 227614 220294 227682 220350
rect 227738 220294 258278 220350
rect 258334 220294 258402 220350
rect 258458 220294 288998 220350
rect 289054 220294 289122 220350
rect 289178 220294 319718 220350
rect 319774 220294 319842 220350
rect 319898 220294 350438 220350
rect 350494 220294 350562 220350
rect 350618 220294 381158 220350
rect 381214 220294 381282 220350
rect 381338 220294 411878 220350
rect 411934 220294 412002 220350
rect 412058 220294 442598 220350
rect 442654 220294 442722 220350
rect 442778 220294 473318 220350
rect 473374 220294 473442 220350
rect 473498 220294 504038 220350
rect 504094 220294 504162 220350
rect 504218 220294 534758 220350
rect 534814 220294 534882 220350
rect 534938 220294 565478 220350
rect 565534 220294 565602 220350
rect 565658 220294 589194 220350
rect 589250 220294 589318 220350
rect 589374 220294 589442 220350
rect 589498 220294 589566 220350
rect 589622 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597980 220350
rect -1916 220226 597980 220294
rect -1916 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 5514 220226
rect 5570 220170 5638 220226
rect 5694 220170 5762 220226
rect 5818 220170 5886 220226
rect 5942 220170 12518 220226
rect 12574 220170 12642 220226
rect 12698 220170 43238 220226
rect 43294 220170 43362 220226
rect 43418 220170 73958 220226
rect 74014 220170 74082 220226
rect 74138 220170 104678 220226
rect 104734 220170 104802 220226
rect 104858 220170 135398 220226
rect 135454 220170 135522 220226
rect 135578 220170 166118 220226
rect 166174 220170 166242 220226
rect 166298 220170 196838 220226
rect 196894 220170 196962 220226
rect 197018 220170 227558 220226
rect 227614 220170 227682 220226
rect 227738 220170 258278 220226
rect 258334 220170 258402 220226
rect 258458 220170 288998 220226
rect 289054 220170 289122 220226
rect 289178 220170 319718 220226
rect 319774 220170 319842 220226
rect 319898 220170 350438 220226
rect 350494 220170 350562 220226
rect 350618 220170 381158 220226
rect 381214 220170 381282 220226
rect 381338 220170 411878 220226
rect 411934 220170 412002 220226
rect 412058 220170 442598 220226
rect 442654 220170 442722 220226
rect 442778 220170 473318 220226
rect 473374 220170 473442 220226
rect 473498 220170 504038 220226
rect 504094 220170 504162 220226
rect 504218 220170 534758 220226
rect 534814 220170 534882 220226
rect 534938 220170 565478 220226
rect 565534 220170 565602 220226
rect 565658 220170 589194 220226
rect 589250 220170 589318 220226
rect 589374 220170 589442 220226
rect 589498 220170 589566 220226
rect 589622 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597980 220226
rect -1916 220102 597980 220170
rect -1916 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 5514 220102
rect 5570 220046 5638 220102
rect 5694 220046 5762 220102
rect 5818 220046 5886 220102
rect 5942 220046 12518 220102
rect 12574 220046 12642 220102
rect 12698 220046 43238 220102
rect 43294 220046 43362 220102
rect 43418 220046 73958 220102
rect 74014 220046 74082 220102
rect 74138 220046 104678 220102
rect 104734 220046 104802 220102
rect 104858 220046 135398 220102
rect 135454 220046 135522 220102
rect 135578 220046 166118 220102
rect 166174 220046 166242 220102
rect 166298 220046 196838 220102
rect 196894 220046 196962 220102
rect 197018 220046 227558 220102
rect 227614 220046 227682 220102
rect 227738 220046 258278 220102
rect 258334 220046 258402 220102
rect 258458 220046 288998 220102
rect 289054 220046 289122 220102
rect 289178 220046 319718 220102
rect 319774 220046 319842 220102
rect 319898 220046 350438 220102
rect 350494 220046 350562 220102
rect 350618 220046 381158 220102
rect 381214 220046 381282 220102
rect 381338 220046 411878 220102
rect 411934 220046 412002 220102
rect 412058 220046 442598 220102
rect 442654 220046 442722 220102
rect 442778 220046 473318 220102
rect 473374 220046 473442 220102
rect 473498 220046 504038 220102
rect 504094 220046 504162 220102
rect 504218 220046 534758 220102
rect 534814 220046 534882 220102
rect 534938 220046 565478 220102
rect 565534 220046 565602 220102
rect 565658 220046 589194 220102
rect 589250 220046 589318 220102
rect 589374 220046 589442 220102
rect 589498 220046 589566 220102
rect 589622 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597980 220102
rect -1916 219978 597980 220046
rect -1916 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 5514 219978
rect 5570 219922 5638 219978
rect 5694 219922 5762 219978
rect 5818 219922 5886 219978
rect 5942 219922 12518 219978
rect 12574 219922 12642 219978
rect 12698 219922 43238 219978
rect 43294 219922 43362 219978
rect 43418 219922 73958 219978
rect 74014 219922 74082 219978
rect 74138 219922 104678 219978
rect 104734 219922 104802 219978
rect 104858 219922 135398 219978
rect 135454 219922 135522 219978
rect 135578 219922 166118 219978
rect 166174 219922 166242 219978
rect 166298 219922 196838 219978
rect 196894 219922 196962 219978
rect 197018 219922 227558 219978
rect 227614 219922 227682 219978
rect 227738 219922 258278 219978
rect 258334 219922 258402 219978
rect 258458 219922 288998 219978
rect 289054 219922 289122 219978
rect 289178 219922 319718 219978
rect 319774 219922 319842 219978
rect 319898 219922 350438 219978
rect 350494 219922 350562 219978
rect 350618 219922 381158 219978
rect 381214 219922 381282 219978
rect 381338 219922 411878 219978
rect 411934 219922 412002 219978
rect 412058 219922 442598 219978
rect 442654 219922 442722 219978
rect 442778 219922 473318 219978
rect 473374 219922 473442 219978
rect 473498 219922 504038 219978
rect 504094 219922 504162 219978
rect 504218 219922 534758 219978
rect 534814 219922 534882 219978
rect 534938 219922 565478 219978
rect 565534 219922 565602 219978
rect 565658 219922 589194 219978
rect 589250 219922 589318 219978
rect 589374 219922 589442 219978
rect 589498 219922 589566 219978
rect 589622 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597980 219978
rect -1916 219826 597980 219922
rect -1916 208350 597980 208446
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 27878 208350
rect 27934 208294 28002 208350
rect 28058 208294 58598 208350
rect 58654 208294 58722 208350
rect 58778 208294 89318 208350
rect 89374 208294 89442 208350
rect 89498 208294 120038 208350
rect 120094 208294 120162 208350
rect 120218 208294 150758 208350
rect 150814 208294 150882 208350
rect 150938 208294 181478 208350
rect 181534 208294 181602 208350
rect 181658 208294 212198 208350
rect 212254 208294 212322 208350
rect 212378 208294 242918 208350
rect 242974 208294 243042 208350
rect 243098 208294 273638 208350
rect 273694 208294 273762 208350
rect 273818 208294 304358 208350
rect 304414 208294 304482 208350
rect 304538 208294 335078 208350
rect 335134 208294 335202 208350
rect 335258 208294 365798 208350
rect 365854 208294 365922 208350
rect 365978 208294 396518 208350
rect 396574 208294 396642 208350
rect 396698 208294 427238 208350
rect 427294 208294 427362 208350
rect 427418 208294 457958 208350
rect 458014 208294 458082 208350
rect 458138 208294 488678 208350
rect 488734 208294 488802 208350
rect 488858 208294 519398 208350
rect 519454 208294 519522 208350
rect 519578 208294 550118 208350
rect 550174 208294 550242 208350
rect 550298 208294 592914 208350
rect 592970 208294 593038 208350
rect 593094 208294 593162 208350
rect 593218 208294 593286 208350
rect 593342 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect -1916 208226 597980 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 27878 208226
rect 27934 208170 28002 208226
rect 28058 208170 58598 208226
rect 58654 208170 58722 208226
rect 58778 208170 89318 208226
rect 89374 208170 89442 208226
rect 89498 208170 120038 208226
rect 120094 208170 120162 208226
rect 120218 208170 150758 208226
rect 150814 208170 150882 208226
rect 150938 208170 181478 208226
rect 181534 208170 181602 208226
rect 181658 208170 212198 208226
rect 212254 208170 212322 208226
rect 212378 208170 242918 208226
rect 242974 208170 243042 208226
rect 243098 208170 273638 208226
rect 273694 208170 273762 208226
rect 273818 208170 304358 208226
rect 304414 208170 304482 208226
rect 304538 208170 335078 208226
rect 335134 208170 335202 208226
rect 335258 208170 365798 208226
rect 365854 208170 365922 208226
rect 365978 208170 396518 208226
rect 396574 208170 396642 208226
rect 396698 208170 427238 208226
rect 427294 208170 427362 208226
rect 427418 208170 457958 208226
rect 458014 208170 458082 208226
rect 458138 208170 488678 208226
rect 488734 208170 488802 208226
rect 488858 208170 519398 208226
rect 519454 208170 519522 208226
rect 519578 208170 550118 208226
rect 550174 208170 550242 208226
rect 550298 208170 592914 208226
rect 592970 208170 593038 208226
rect 593094 208170 593162 208226
rect 593218 208170 593286 208226
rect 593342 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect -1916 208102 597980 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 27878 208102
rect 27934 208046 28002 208102
rect 28058 208046 58598 208102
rect 58654 208046 58722 208102
rect 58778 208046 89318 208102
rect 89374 208046 89442 208102
rect 89498 208046 120038 208102
rect 120094 208046 120162 208102
rect 120218 208046 150758 208102
rect 150814 208046 150882 208102
rect 150938 208046 181478 208102
rect 181534 208046 181602 208102
rect 181658 208046 212198 208102
rect 212254 208046 212322 208102
rect 212378 208046 242918 208102
rect 242974 208046 243042 208102
rect 243098 208046 273638 208102
rect 273694 208046 273762 208102
rect 273818 208046 304358 208102
rect 304414 208046 304482 208102
rect 304538 208046 335078 208102
rect 335134 208046 335202 208102
rect 335258 208046 365798 208102
rect 365854 208046 365922 208102
rect 365978 208046 396518 208102
rect 396574 208046 396642 208102
rect 396698 208046 427238 208102
rect 427294 208046 427362 208102
rect 427418 208046 457958 208102
rect 458014 208046 458082 208102
rect 458138 208046 488678 208102
rect 488734 208046 488802 208102
rect 488858 208046 519398 208102
rect 519454 208046 519522 208102
rect 519578 208046 550118 208102
rect 550174 208046 550242 208102
rect 550298 208046 592914 208102
rect 592970 208046 593038 208102
rect 593094 208046 593162 208102
rect 593218 208046 593286 208102
rect 593342 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect -1916 207978 597980 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 27878 207978
rect 27934 207922 28002 207978
rect 28058 207922 58598 207978
rect 58654 207922 58722 207978
rect 58778 207922 89318 207978
rect 89374 207922 89442 207978
rect 89498 207922 120038 207978
rect 120094 207922 120162 207978
rect 120218 207922 150758 207978
rect 150814 207922 150882 207978
rect 150938 207922 181478 207978
rect 181534 207922 181602 207978
rect 181658 207922 212198 207978
rect 212254 207922 212322 207978
rect 212378 207922 242918 207978
rect 242974 207922 243042 207978
rect 243098 207922 273638 207978
rect 273694 207922 273762 207978
rect 273818 207922 304358 207978
rect 304414 207922 304482 207978
rect 304538 207922 335078 207978
rect 335134 207922 335202 207978
rect 335258 207922 365798 207978
rect 365854 207922 365922 207978
rect 365978 207922 396518 207978
rect 396574 207922 396642 207978
rect 396698 207922 427238 207978
rect 427294 207922 427362 207978
rect 427418 207922 457958 207978
rect 458014 207922 458082 207978
rect 458138 207922 488678 207978
rect 488734 207922 488802 207978
rect 488858 207922 519398 207978
rect 519454 207922 519522 207978
rect 519578 207922 550118 207978
rect 550174 207922 550242 207978
rect 550298 207922 592914 207978
rect 592970 207922 593038 207978
rect 593094 207922 593162 207978
rect 593218 207922 593286 207978
rect 593342 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect -1916 207826 597980 207922
rect -1916 202350 597980 202446
rect -1916 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 5514 202350
rect 5570 202294 5638 202350
rect 5694 202294 5762 202350
rect 5818 202294 5886 202350
rect 5942 202294 12518 202350
rect 12574 202294 12642 202350
rect 12698 202294 43238 202350
rect 43294 202294 43362 202350
rect 43418 202294 73958 202350
rect 74014 202294 74082 202350
rect 74138 202294 104678 202350
rect 104734 202294 104802 202350
rect 104858 202294 135398 202350
rect 135454 202294 135522 202350
rect 135578 202294 166118 202350
rect 166174 202294 166242 202350
rect 166298 202294 196838 202350
rect 196894 202294 196962 202350
rect 197018 202294 227558 202350
rect 227614 202294 227682 202350
rect 227738 202294 258278 202350
rect 258334 202294 258402 202350
rect 258458 202294 288998 202350
rect 289054 202294 289122 202350
rect 289178 202294 319718 202350
rect 319774 202294 319842 202350
rect 319898 202294 350438 202350
rect 350494 202294 350562 202350
rect 350618 202294 381158 202350
rect 381214 202294 381282 202350
rect 381338 202294 411878 202350
rect 411934 202294 412002 202350
rect 412058 202294 442598 202350
rect 442654 202294 442722 202350
rect 442778 202294 473318 202350
rect 473374 202294 473442 202350
rect 473498 202294 504038 202350
rect 504094 202294 504162 202350
rect 504218 202294 534758 202350
rect 534814 202294 534882 202350
rect 534938 202294 565478 202350
rect 565534 202294 565602 202350
rect 565658 202294 589194 202350
rect 589250 202294 589318 202350
rect 589374 202294 589442 202350
rect 589498 202294 589566 202350
rect 589622 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597980 202350
rect -1916 202226 597980 202294
rect -1916 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 5514 202226
rect 5570 202170 5638 202226
rect 5694 202170 5762 202226
rect 5818 202170 5886 202226
rect 5942 202170 12518 202226
rect 12574 202170 12642 202226
rect 12698 202170 43238 202226
rect 43294 202170 43362 202226
rect 43418 202170 73958 202226
rect 74014 202170 74082 202226
rect 74138 202170 104678 202226
rect 104734 202170 104802 202226
rect 104858 202170 135398 202226
rect 135454 202170 135522 202226
rect 135578 202170 166118 202226
rect 166174 202170 166242 202226
rect 166298 202170 196838 202226
rect 196894 202170 196962 202226
rect 197018 202170 227558 202226
rect 227614 202170 227682 202226
rect 227738 202170 258278 202226
rect 258334 202170 258402 202226
rect 258458 202170 288998 202226
rect 289054 202170 289122 202226
rect 289178 202170 319718 202226
rect 319774 202170 319842 202226
rect 319898 202170 350438 202226
rect 350494 202170 350562 202226
rect 350618 202170 381158 202226
rect 381214 202170 381282 202226
rect 381338 202170 411878 202226
rect 411934 202170 412002 202226
rect 412058 202170 442598 202226
rect 442654 202170 442722 202226
rect 442778 202170 473318 202226
rect 473374 202170 473442 202226
rect 473498 202170 504038 202226
rect 504094 202170 504162 202226
rect 504218 202170 534758 202226
rect 534814 202170 534882 202226
rect 534938 202170 565478 202226
rect 565534 202170 565602 202226
rect 565658 202170 589194 202226
rect 589250 202170 589318 202226
rect 589374 202170 589442 202226
rect 589498 202170 589566 202226
rect 589622 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597980 202226
rect -1916 202102 597980 202170
rect -1916 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 5514 202102
rect 5570 202046 5638 202102
rect 5694 202046 5762 202102
rect 5818 202046 5886 202102
rect 5942 202046 12518 202102
rect 12574 202046 12642 202102
rect 12698 202046 43238 202102
rect 43294 202046 43362 202102
rect 43418 202046 73958 202102
rect 74014 202046 74082 202102
rect 74138 202046 104678 202102
rect 104734 202046 104802 202102
rect 104858 202046 135398 202102
rect 135454 202046 135522 202102
rect 135578 202046 166118 202102
rect 166174 202046 166242 202102
rect 166298 202046 196838 202102
rect 196894 202046 196962 202102
rect 197018 202046 227558 202102
rect 227614 202046 227682 202102
rect 227738 202046 258278 202102
rect 258334 202046 258402 202102
rect 258458 202046 288998 202102
rect 289054 202046 289122 202102
rect 289178 202046 319718 202102
rect 319774 202046 319842 202102
rect 319898 202046 350438 202102
rect 350494 202046 350562 202102
rect 350618 202046 381158 202102
rect 381214 202046 381282 202102
rect 381338 202046 411878 202102
rect 411934 202046 412002 202102
rect 412058 202046 442598 202102
rect 442654 202046 442722 202102
rect 442778 202046 473318 202102
rect 473374 202046 473442 202102
rect 473498 202046 504038 202102
rect 504094 202046 504162 202102
rect 504218 202046 534758 202102
rect 534814 202046 534882 202102
rect 534938 202046 565478 202102
rect 565534 202046 565602 202102
rect 565658 202046 589194 202102
rect 589250 202046 589318 202102
rect 589374 202046 589442 202102
rect 589498 202046 589566 202102
rect 589622 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597980 202102
rect -1916 201978 597980 202046
rect -1916 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 5514 201978
rect 5570 201922 5638 201978
rect 5694 201922 5762 201978
rect 5818 201922 5886 201978
rect 5942 201922 12518 201978
rect 12574 201922 12642 201978
rect 12698 201922 43238 201978
rect 43294 201922 43362 201978
rect 43418 201922 73958 201978
rect 74014 201922 74082 201978
rect 74138 201922 104678 201978
rect 104734 201922 104802 201978
rect 104858 201922 135398 201978
rect 135454 201922 135522 201978
rect 135578 201922 166118 201978
rect 166174 201922 166242 201978
rect 166298 201922 196838 201978
rect 196894 201922 196962 201978
rect 197018 201922 227558 201978
rect 227614 201922 227682 201978
rect 227738 201922 258278 201978
rect 258334 201922 258402 201978
rect 258458 201922 288998 201978
rect 289054 201922 289122 201978
rect 289178 201922 319718 201978
rect 319774 201922 319842 201978
rect 319898 201922 350438 201978
rect 350494 201922 350562 201978
rect 350618 201922 381158 201978
rect 381214 201922 381282 201978
rect 381338 201922 411878 201978
rect 411934 201922 412002 201978
rect 412058 201922 442598 201978
rect 442654 201922 442722 201978
rect 442778 201922 473318 201978
rect 473374 201922 473442 201978
rect 473498 201922 504038 201978
rect 504094 201922 504162 201978
rect 504218 201922 534758 201978
rect 534814 201922 534882 201978
rect 534938 201922 565478 201978
rect 565534 201922 565602 201978
rect 565658 201922 589194 201978
rect 589250 201922 589318 201978
rect 589374 201922 589442 201978
rect 589498 201922 589566 201978
rect 589622 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597980 201978
rect -1916 201826 597980 201922
rect -1916 190350 597980 190446
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 27878 190350
rect 27934 190294 28002 190350
rect 28058 190294 58598 190350
rect 58654 190294 58722 190350
rect 58778 190294 89318 190350
rect 89374 190294 89442 190350
rect 89498 190294 120038 190350
rect 120094 190294 120162 190350
rect 120218 190294 150758 190350
rect 150814 190294 150882 190350
rect 150938 190294 181478 190350
rect 181534 190294 181602 190350
rect 181658 190294 212198 190350
rect 212254 190294 212322 190350
rect 212378 190294 242918 190350
rect 242974 190294 243042 190350
rect 243098 190294 273638 190350
rect 273694 190294 273762 190350
rect 273818 190294 304358 190350
rect 304414 190294 304482 190350
rect 304538 190294 335078 190350
rect 335134 190294 335202 190350
rect 335258 190294 365798 190350
rect 365854 190294 365922 190350
rect 365978 190294 396518 190350
rect 396574 190294 396642 190350
rect 396698 190294 427238 190350
rect 427294 190294 427362 190350
rect 427418 190294 457958 190350
rect 458014 190294 458082 190350
rect 458138 190294 488678 190350
rect 488734 190294 488802 190350
rect 488858 190294 519398 190350
rect 519454 190294 519522 190350
rect 519578 190294 550118 190350
rect 550174 190294 550242 190350
rect 550298 190294 592914 190350
rect 592970 190294 593038 190350
rect 593094 190294 593162 190350
rect 593218 190294 593286 190350
rect 593342 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect -1916 190226 597980 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 27878 190226
rect 27934 190170 28002 190226
rect 28058 190170 58598 190226
rect 58654 190170 58722 190226
rect 58778 190170 89318 190226
rect 89374 190170 89442 190226
rect 89498 190170 120038 190226
rect 120094 190170 120162 190226
rect 120218 190170 150758 190226
rect 150814 190170 150882 190226
rect 150938 190170 181478 190226
rect 181534 190170 181602 190226
rect 181658 190170 212198 190226
rect 212254 190170 212322 190226
rect 212378 190170 242918 190226
rect 242974 190170 243042 190226
rect 243098 190170 273638 190226
rect 273694 190170 273762 190226
rect 273818 190170 304358 190226
rect 304414 190170 304482 190226
rect 304538 190170 335078 190226
rect 335134 190170 335202 190226
rect 335258 190170 365798 190226
rect 365854 190170 365922 190226
rect 365978 190170 396518 190226
rect 396574 190170 396642 190226
rect 396698 190170 427238 190226
rect 427294 190170 427362 190226
rect 427418 190170 457958 190226
rect 458014 190170 458082 190226
rect 458138 190170 488678 190226
rect 488734 190170 488802 190226
rect 488858 190170 519398 190226
rect 519454 190170 519522 190226
rect 519578 190170 550118 190226
rect 550174 190170 550242 190226
rect 550298 190170 592914 190226
rect 592970 190170 593038 190226
rect 593094 190170 593162 190226
rect 593218 190170 593286 190226
rect 593342 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect -1916 190102 597980 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 27878 190102
rect 27934 190046 28002 190102
rect 28058 190046 58598 190102
rect 58654 190046 58722 190102
rect 58778 190046 89318 190102
rect 89374 190046 89442 190102
rect 89498 190046 120038 190102
rect 120094 190046 120162 190102
rect 120218 190046 150758 190102
rect 150814 190046 150882 190102
rect 150938 190046 181478 190102
rect 181534 190046 181602 190102
rect 181658 190046 212198 190102
rect 212254 190046 212322 190102
rect 212378 190046 242918 190102
rect 242974 190046 243042 190102
rect 243098 190046 273638 190102
rect 273694 190046 273762 190102
rect 273818 190046 304358 190102
rect 304414 190046 304482 190102
rect 304538 190046 335078 190102
rect 335134 190046 335202 190102
rect 335258 190046 365798 190102
rect 365854 190046 365922 190102
rect 365978 190046 396518 190102
rect 396574 190046 396642 190102
rect 396698 190046 427238 190102
rect 427294 190046 427362 190102
rect 427418 190046 457958 190102
rect 458014 190046 458082 190102
rect 458138 190046 488678 190102
rect 488734 190046 488802 190102
rect 488858 190046 519398 190102
rect 519454 190046 519522 190102
rect 519578 190046 550118 190102
rect 550174 190046 550242 190102
rect 550298 190046 592914 190102
rect 592970 190046 593038 190102
rect 593094 190046 593162 190102
rect 593218 190046 593286 190102
rect 593342 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect -1916 189978 597980 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 27878 189978
rect 27934 189922 28002 189978
rect 28058 189922 58598 189978
rect 58654 189922 58722 189978
rect 58778 189922 89318 189978
rect 89374 189922 89442 189978
rect 89498 189922 120038 189978
rect 120094 189922 120162 189978
rect 120218 189922 150758 189978
rect 150814 189922 150882 189978
rect 150938 189922 181478 189978
rect 181534 189922 181602 189978
rect 181658 189922 212198 189978
rect 212254 189922 212322 189978
rect 212378 189922 242918 189978
rect 242974 189922 243042 189978
rect 243098 189922 273638 189978
rect 273694 189922 273762 189978
rect 273818 189922 304358 189978
rect 304414 189922 304482 189978
rect 304538 189922 335078 189978
rect 335134 189922 335202 189978
rect 335258 189922 365798 189978
rect 365854 189922 365922 189978
rect 365978 189922 396518 189978
rect 396574 189922 396642 189978
rect 396698 189922 427238 189978
rect 427294 189922 427362 189978
rect 427418 189922 457958 189978
rect 458014 189922 458082 189978
rect 458138 189922 488678 189978
rect 488734 189922 488802 189978
rect 488858 189922 519398 189978
rect 519454 189922 519522 189978
rect 519578 189922 550118 189978
rect 550174 189922 550242 189978
rect 550298 189922 592914 189978
rect 592970 189922 593038 189978
rect 593094 189922 593162 189978
rect 593218 189922 593286 189978
rect 593342 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect -1916 189826 597980 189922
rect -1916 184350 597980 184446
rect -1916 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 5514 184350
rect 5570 184294 5638 184350
rect 5694 184294 5762 184350
rect 5818 184294 5886 184350
rect 5942 184294 12518 184350
rect 12574 184294 12642 184350
rect 12698 184294 43238 184350
rect 43294 184294 43362 184350
rect 43418 184294 73958 184350
rect 74014 184294 74082 184350
rect 74138 184294 104678 184350
rect 104734 184294 104802 184350
rect 104858 184294 135398 184350
rect 135454 184294 135522 184350
rect 135578 184294 166118 184350
rect 166174 184294 166242 184350
rect 166298 184294 196838 184350
rect 196894 184294 196962 184350
rect 197018 184294 227558 184350
rect 227614 184294 227682 184350
rect 227738 184294 258278 184350
rect 258334 184294 258402 184350
rect 258458 184294 288998 184350
rect 289054 184294 289122 184350
rect 289178 184294 319718 184350
rect 319774 184294 319842 184350
rect 319898 184294 350438 184350
rect 350494 184294 350562 184350
rect 350618 184294 381158 184350
rect 381214 184294 381282 184350
rect 381338 184294 411878 184350
rect 411934 184294 412002 184350
rect 412058 184294 442598 184350
rect 442654 184294 442722 184350
rect 442778 184294 473318 184350
rect 473374 184294 473442 184350
rect 473498 184294 504038 184350
rect 504094 184294 504162 184350
rect 504218 184294 534758 184350
rect 534814 184294 534882 184350
rect 534938 184294 565478 184350
rect 565534 184294 565602 184350
rect 565658 184294 589194 184350
rect 589250 184294 589318 184350
rect 589374 184294 589442 184350
rect 589498 184294 589566 184350
rect 589622 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597980 184350
rect -1916 184226 597980 184294
rect -1916 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 5514 184226
rect 5570 184170 5638 184226
rect 5694 184170 5762 184226
rect 5818 184170 5886 184226
rect 5942 184170 12518 184226
rect 12574 184170 12642 184226
rect 12698 184170 43238 184226
rect 43294 184170 43362 184226
rect 43418 184170 73958 184226
rect 74014 184170 74082 184226
rect 74138 184170 104678 184226
rect 104734 184170 104802 184226
rect 104858 184170 135398 184226
rect 135454 184170 135522 184226
rect 135578 184170 166118 184226
rect 166174 184170 166242 184226
rect 166298 184170 196838 184226
rect 196894 184170 196962 184226
rect 197018 184170 227558 184226
rect 227614 184170 227682 184226
rect 227738 184170 258278 184226
rect 258334 184170 258402 184226
rect 258458 184170 288998 184226
rect 289054 184170 289122 184226
rect 289178 184170 319718 184226
rect 319774 184170 319842 184226
rect 319898 184170 350438 184226
rect 350494 184170 350562 184226
rect 350618 184170 381158 184226
rect 381214 184170 381282 184226
rect 381338 184170 411878 184226
rect 411934 184170 412002 184226
rect 412058 184170 442598 184226
rect 442654 184170 442722 184226
rect 442778 184170 473318 184226
rect 473374 184170 473442 184226
rect 473498 184170 504038 184226
rect 504094 184170 504162 184226
rect 504218 184170 534758 184226
rect 534814 184170 534882 184226
rect 534938 184170 565478 184226
rect 565534 184170 565602 184226
rect 565658 184170 589194 184226
rect 589250 184170 589318 184226
rect 589374 184170 589442 184226
rect 589498 184170 589566 184226
rect 589622 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597980 184226
rect -1916 184102 597980 184170
rect -1916 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 5514 184102
rect 5570 184046 5638 184102
rect 5694 184046 5762 184102
rect 5818 184046 5886 184102
rect 5942 184046 12518 184102
rect 12574 184046 12642 184102
rect 12698 184046 43238 184102
rect 43294 184046 43362 184102
rect 43418 184046 73958 184102
rect 74014 184046 74082 184102
rect 74138 184046 104678 184102
rect 104734 184046 104802 184102
rect 104858 184046 135398 184102
rect 135454 184046 135522 184102
rect 135578 184046 166118 184102
rect 166174 184046 166242 184102
rect 166298 184046 196838 184102
rect 196894 184046 196962 184102
rect 197018 184046 227558 184102
rect 227614 184046 227682 184102
rect 227738 184046 258278 184102
rect 258334 184046 258402 184102
rect 258458 184046 288998 184102
rect 289054 184046 289122 184102
rect 289178 184046 319718 184102
rect 319774 184046 319842 184102
rect 319898 184046 350438 184102
rect 350494 184046 350562 184102
rect 350618 184046 381158 184102
rect 381214 184046 381282 184102
rect 381338 184046 411878 184102
rect 411934 184046 412002 184102
rect 412058 184046 442598 184102
rect 442654 184046 442722 184102
rect 442778 184046 473318 184102
rect 473374 184046 473442 184102
rect 473498 184046 504038 184102
rect 504094 184046 504162 184102
rect 504218 184046 534758 184102
rect 534814 184046 534882 184102
rect 534938 184046 565478 184102
rect 565534 184046 565602 184102
rect 565658 184046 589194 184102
rect 589250 184046 589318 184102
rect 589374 184046 589442 184102
rect 589498 184046 589566 184102
rect 589622 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597980 184102
rect -1916 183978 597980 184046
rect -1916 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 5514 183978
rect 5570 183922 5638 183978
rect 5694 183922 5762 183978
rect 5818 183922 5886 183978
rect 5942 183922 12518 183978
rect 12574 183922 12642 183978
rect 12698 183922 43238 183978
rect 43294 183922 43362 183978
rect 43418 183922 73958 183978
rect 74014 183922 74082 183978
rect 74138 183922 104678 183978
rect 104734 183922 104802 183978
rect 104858 183922 135398 183978
rect 135454 183922 135522 183978
rect 135578 183922 166118 183978
rect 166174 183922 166242 183978
rect 166298 183922 196838 183978
rect 196894 183922 196962 183978
rect 197018 183922 227558 183978
rect 227614 183922 227682 183978
rect 227738 183922 258278 183978
rect 258334 183922 258402 183978
rect 258458 183922 288998 183978
rect 289054 183922 289122 183978
rect 289178 183922 319718 183978
rect 319774 183922 319842 183978
rect 319898 183922 350438 183978
rect 350494 183922 350562 183978
rect 350618 183922 381158 183978
rect 381214 183922 381282 183978
rect 381338 183922 411878 183978
rect 411934 183922 412002 183978
rect 412058 183922 442598 183978
rect 442654 183922 442722 183978
rect 442778 183922 473318 183978
rect 473374 183922 473442 183978
rect 473498 183922 504038 183978
rect 504094 183922 504162 183978
rect 504218 183922 534758 183978
rect 534814 183922 534882 183978
rect 534938 183922 565478 183978
rect 565534 183922 565602 183978
rect 565658 183922 589194 183978
rect 589250 183922 589318 183978
rect 589374 183922 589442 183978
rect 589498 183922 589566 183978
rect 589622 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597980 183978
rect -1916 183826 597980 183922
rect -1916 172350 597980 172446
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 27878 172350
rect 27934 172294 28002 172350
rect 28058 172294 58598 172350
rect 58654 172294 58722 172350
rect 58778 172294 89318 172350
rect 89374 172294 89442 172350
rect 89498 172294 120038 172350
rect 120094 172294 120162 172350
rect 120218 172294 150758 172350
rect 150814 172294 150882 172350
rect 150938 172294 181478 172350
rect 181534 172294 181602 172350
rect 181658 172294 212198 172350
rect 212254 172294 212322 172350
rect 212378 172294 242918 172350
rect 242974 172294 243042 172350
rect 243098 172294 273638 172350
rect 273694 172294 273762 172350
rect 273818 172294 304358 172350
rect 304414 172294 304482 172350
rect 304538 172294 335078 172350
rect 335134 172294 335202 172350
rect 335258 172294 365798 172350
rect 365854 172294 365922 172350
rect 365978 172294 396518 172350
rect 396574 172294 396642 172350
rect 396698 172294 427238 172350
rect 427294 172294 427362 172350
rect 427418 172294 457958 172350
rect 458014 172294 458082 172350
rect 458138 172294 488678 172350
rect 488734 172294 488802 172350
rect 488858 172294 519398 172350
rect 519454 172294 519522 172350
rect 519578 172294 550118 172350
rect 550174 172294 550242 172350
rect 550298 172294 592914 172350
rect 592970 172294 593038 172350
rect 593094 172294 593162 172350
rect 593218 172294 593286 172350
rect 593342 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect -1916 172226 597980 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 27878 172226
rect 27934 172170 28002 172226
rect 28058 172170 58598 172226
rect 58654 172170 58722 172226
rect 58778 172170 89318 172226
rect 89374 172170 89442 172226
rect 89498 172170 120038 172226
rect 120094 172170 120162 172226
rect 120218 172170 150758 172226
rect 150814 172170 150882 172226
rect 150938 172170 181478 172226
rect 181534 172170 181602 172226
rect 181658 172170 212198 172226
rect 212254 172170 212322 172226
rect 212378 172170 242918 172226
rect 242974 172170 243042 172226
rect 243098 172170 273638 172226
rect 273694 172170 273762 172226
rect 273818 172170 304358 172226
rect 304414 172170 304482 172226
rect 304538 172170 335078 172226
rect 335134 172170 335202 172226
rect 335258 172170 365798 172226
rect 365854 172170 365922 172226
rect 365978 172170 396518 172226
rect 396574 172170 396642 172226
rect 396698 172170 427238 172226
rect 427294 172170 427362 172226
rect 427418 172170 457958 172226
rect 458014 172170 458082 172226
rect 458138 172170 488678 172226
rect 488734 172170 488802 172226
rect 488858 172170 519398 172226
rect 519454 172170 519522 172226
rect 519578 172170 550118 172226
rect 550174 172170 550242 172226
rect 550298 172170 592914 172226
rect 592970 172170 593038 172226
rect 593094 172170 593162 172226
rect 593218 172170 593286 172226
rect 593342 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect -1916 172102 597980 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 27878 172102
rect 27934 172046 28002 172102
rect 28058 172046 58598 172102
rect 58654 172046 58722 172102
rect 58778 172046 89318 172102
rect 89374 172046 89442 172102
rect 89498 172046 120038 172102
rect 120094 172046 120162 172102
rect 120218 172046 150758 172102
rect 150814 172046 150882 172102
rect 150938 172046 181478 172102
rect 181534 172046 181602 172102
rect 181658 172046 212198 172102
rect 212254 172046 212322 172102
rect 212378 172046 242918 172102
rect 242974 172046 243042 172102
rect 243098 172046 273638 172102
rect 273694 172046 273762 172102
rect 273818 172046 304358 172102
rect 304414 172046 304482 172102
rect 304538 172046 335078 172102
rect 335134 172046 335202 172102
rect 335258 172046 365798 172102
rect 365854 172046 365922 172102
rect 365978 172046 396518 172102
rect 396574 172046 396642 172102
rect 396698 172046 427238 172102
rect 427294 172046 427362 172102
rect 427418 172046 457958 172102
rect 458014 172046 458082 172102
rect 458138 172046 488678 172102
rect 488734 172046 488802 172102
rect 488858 172046 519398 172102
rect 519454 172046 519522 172102
rect 519578 172046 550118 172102
rect 550174 172046 550242 172102
rect 550298 172046 592914 172102
rect 592970 172046 593038 172102
rect 593094 172046 593162 172102
rect 593218 172046 593286 172102
rect 593342 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect -1916 171978 597980 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 27878 171978
rect 27934 171922 28002 171978
rect 28058 171922 58598 171978
rect 58654 171922 58722 171978
rect 58778 171922 89318 171978
rect 89374 171922 89442 171978
rect 89498 171922 120038 171978
rect 120094 171922 120162 171978
rect 120218 171922 150758 171978
rect 150814 171922 150882 171978
rect 150938 171922 181478 171978
rect 181534 171922 181602 171978
rect 181658 171922 212198 171978
rect 212254 171922 212322 171978
rect 212378 171922 242918 171978
rect 242974 171922 243042 171978
rect 243098 171922 273638 171978
rect 273694 171922 273762 171978
rect 273818 171922 304358 171978
rect 304414 171922 304482 171978
rect 304538 171922 335078 171978
rect 335134 171922 335202 171978
rect 335258 171922 365798 171978
rect 365854 171922 365922 171978
rect 365978 171922 396518 171978
rect 396574 171922 396642 171978
rect 396698 171922 427238 171978
rect 427294 171922 427362 171978
rect 427418 171922 457958 171978
rect 458014 171922 458082 171978
rect 458138 171922 488678 171978
rect 488734 171922 488802 171978
rect 488858 171922 519398 171978
rect 519454 171922 519522 171978
rect 519578 171922 550118 171978
rect 550174 171922 550242 171978
rect 550298 171922 592914 171978
rect 592970 171922 593038 171978
rect 593094 171922 593162 171978
rect 593218 171922 593286 171978
rect 593342 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect -1916 171826 597980 171922
rect -1916 166350 597980 166446
rect -1916 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 5514 166350
rect 5570 166294 5638 166350
rect 5694 166294 5762 166350
rect 5818 166294 5886 166350
rect 5942 166294 12518 166350
rect 12574 166294 12642 166350
rect 12698 166294 43238 166350
rect 43294 166294 43362 166350
rect 43418 166294 73958 166350
rect 74014 166294 74082 166350
rect 74138 166294 104678 166350
rect 104734 166294 104802 166350
rect 104858 166294 135398 166350
rect 135454 166294 135522 166350
rect 135578 166294 166118 166350
rect 166174 166294 166242 166350
rect 166298 166294 196838 166350
rect 196894 166294 196962 166350
rect 197018 166294 227558 166350
rect 227614 166294 227682 166350
rect 227738 166294 258278 166350
rect 258334 166294 258402 166350
rect 258458 166294 288998 166350
rect 289054 166294 289122 166350
rect 289178 166294 319718 166350
rect 319774 166294 319842 166350
rect 319898 166294 350438 166350
rect 350494 166294 350562 166350
rect 350618 166294 381158 166350
rect 381214 166294 381282 166350
rect 381338 166294 411878 166350
rect 411934 166294 412002 166350
rect 412058 166294 442598 166350
rect 442654 166294 442722 166350
rect 442778 166294 473318 166350
rect 473374 166294 473442 166350
rect 473498 166294 504038 166350
rect 504094 166294 504162 166350
rect 504218 166294 534758 166350
rect 534814 166294 534882 166350
rect 534938 166294 565478 166350
rect 565534 166294 565602 166350
rect 565658 166294 589194 166350
rect 589250 166294 589318 166350
rect 589374 166294 589442 166350
rect 589498 166294 589566 166350
rect 589622 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597980 166350
rect -1916 166226 597980 166294
rect -1916 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 5514 166226
rect 5570 166170 5638 166226
rect 5694 166170 5762 166226
rect 5818 166170 5886 166226
rect 5942 166170 12518 166226
rect 12574 166170 12642 166226
rect 12698 166170 43238 166226
rect 43294 166170 43362 166226
rect 43418 166170 73958 166226
rect 74014 166170 74082 166226
rect 74138 166170 104678 166226
rect 104734 166170 104802 166226
rect 104858 166170 135398 166226
rect 135454 166170 135522 166226
rect 135578 166170 166118 166226
rect 166174 166170 166242 166226
rect 166298 166170 196838 166226
rect 196894 166170 196962 166226
rect 197018 166170 227558 166226
rect 227614 166170 227682 166226
rect 227738 166170 258278 166226
rect 258334 166170 258402 166226
rect 258458 166170 288998 166226
rect 289054 166170 289122 166226
rect 289178 166170 319718 166226
rect 319774 166170 319842 166226
rect 319898 166170 350438 166226
rect 350494 166170 350562 166226
rect 350618 166170 381158 166226
rect 381214 166170 381282 166226
rect 381338 166170 411878 166226
rect 411934 166170 412002 166226
rect 412058 166170 442598 166226
rect 442654 166170 442722 166226
rect 442778 166170 473318 166226
rect 473374 166170 473442 166226
rect 473498 166170 504038 166226
rect 504094 166170 504162 166226
rect 504218 166170 534758 166226
rect 534814 166170 534882 166226
rect 534938 166170 565478 166226
rect 565534 166170 565602 166226
rect 565658 166170 589194 166226
rect 589250 166170 589318 166226
rect 589374 166170 589442 166226
rect 589498 166170 589566 166226
rect 589622 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597980 166226
rect -1916 166102 597980 166170
rect -1916 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 5514 166102
rect 5570 166046 5638 166102
rect 5694 166046 5762 166102
rect 5818 166046 5886 166102
rect 5942 166046 12518 166102
rect 12574 166046 12642 166102
rect 12698 166046 43238 166102
rect 43294 166046 43362 166102
rect 43418 166046 73958 166102
rect 74014 166046 74082 166102
rect 74138 166046 104678 166102
rect 104734 166046 104802 166102
rect 104858 166046 135398 166102
rect 135454 166046 135522 166102
rect 135578 166046 166118 166102
rect 166174 166046 166242 166102
rect 166298 166046 196838 166102
rect 196894 166046 196962 166102
rect 197018 166046 227558 166102
rect 227614 166046 227682 166102
rect 227738 166046 258278 166102
rect 258334 166046 258402 166102
rect 258458 166046 288998 166102
rect 289054 166046 289122 166102
rect 289178 166046 319718 166102
rect 319774 166046 319842 166102
rect 319898 166046 350438 166102
rect 350494 166046 350562 166102
rect 350618 166046 381158 166102
rect 381214 166046 381282 166102
rect 381338 166046 411878 166102
rect 411934 166046 412002 166102
rect 412058 166046 442598 166102
rect 442654 166046 442722 166102
rect 442778 166046 473318 166102
rect 473374 166046 473442 166102
rect 473498 166046 504038 166102
rect 504094 166046 504162 166102
rect 504218 166046 534758 166102
rect 534814 166046 534882 166102
rect 534938 166046 565478 166102
rect 565534 166046 565602 166102
rect 565658 166046 589194 166102
rect 589250 166046 589318 166102
rect 589374 166046 589442 166102
rect 589498 166046 589566 166102
rect 589622 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597980 166102
rect -1916 165978 597980 166046
rect -1916 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 5514 165978
rect 5570 165922 5638 165978
rect 5694 165922 5762 165978
rect 5818 165922 5886 165978
rect 5942 165922 12518 165978
rect 12574 165922 12642 165978
rect 12698 165922 43238 165978
rect 43294 165922 43362 165978
rect 43418 165922 73958 165978
rect 74014 165922 74082 165978
rect 74138 165922 104678 165978
rect 104734 165922 104802 165978
rect 104858 165922 135398 165978
rect 135454 165922 135522 165978
rect 135578 165922 166118 165978
rect 166174 165922 166242 165978
rect 166298 165922 196838 165978
rect 196894 165922 196962 165978
rect 197018 165922 227558 165978
rect 227614 165922 227682 165978
rect 227738 165922 258278 165978
rect 258334 165922 258402 165978
rect 258458 165922 288998 165978
rect 289054 165922 289122 165978
rect 289178 165922 319718 165978
rect 319774 165922 319842 165978
rect 319898 165922 350438 165978
rect 350494 165922 350562 165978
rect 350618 165922 381158 165978
rect 381214 165922 381282 165978
rect 381338 165922 411878 165978
rect 411934 165922 412002 165978
rect 412058 165922 442598 165978
rect 442654 165922 442722 165978
rect 442778 165922 473318 165978
rect 473374 165922 473442 165978
rect 473498 165922 504038 165978
rect 504094 165922 504162 165978
rect 504218 165922 534758 165978
rect 534814 165922 534882 165978
rect 534938 165922 565478 165978
rect 565534 165922 565602 165978
rect 565658 165922 589194 165978
rect 589250 165922 589318 165978
rect 589374 165922 589442 165978
rect 589498 165922 589566 165978
rect 589622 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597980 165978
rect -1916 165826 597980 165922
rect -1916 154350 597980 154446
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 27878 154350
rect 27934 154294 28002 154350
rect 28058 154294 58598 154350
rect 58654 154294 58722 154350
rect 58778 154294 89318 154350
rect 89374 154294 89442 154350
rect 89498 154294 120038 154350
rect 120094 154294 120162 154350
rect 120218 154294 150758 154350
rect 150814 154294 150882 154350
rect 150938 154294 181478 154350
rect 181534 154294 181602 154350
rect 181658 154294 212198 154350
rect 212254 154294 212322 154350
rect 212378 154294 242918 154350
rect 242974 154294 243042 154350
rect 243098 154294 273638 154350
rect 273694 154294 273762 154350
rect 273818 154294 304358 154350
rect 304414 154294 304482 154350
rect 304538 154294 335078 154350
rect 335134 154294 335202 154350
rect 335258 154294 365798 154350
rect 365854 154294 365922 154350
rect 365978 154294 396518 154350
rect 396574 154294 396642 154350
rect 396698 154294 427238 154350
rect 427294 154294 427362 154350
rect 427418 154294 457958 154350
rect 458014 154294 458082 154350
rect 458138 154294 488678 154350
rect 488734 154294 488802 154350
rect 488858 154294 519398 154350
rect 519454 154294 519522 154350
rect 519578 154294 550118 154350
rect 550174 154294 550242 154350
rect 550298 154294 592914 154350
rect 592970 154294 593038 154350
rect 593094 154294 593162 154350
rect 593218 154294 593286 154350
rect 593342 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect -1916 154226 597980 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 27878 154226
rect 27934 154170 28002 154226
rect 28058 154170 58598 154226
rect 58654 154170 58722 154226
rect 58778 154170 89318 154226
rect 89374 154170 89442 154226
rect 89498 154170 120038 154226
rect 120094 154170 120162 154226
rect 120218 154170 150758 154226
rect 150814 154170 150882 154226
rect 150938 154170 181478 154226
rect 181534 154170 181602 154226
rect 181658 154170 212198 154226
rect 212254 154170 212322 154226
rect 212378 154170 242918 154226
rect 242974 154170 243042 154226
rect 243098 154170 273638 154226
rect 273694 154170 273762 154226
rect 273818 154170 304358 154226
rect 304414 154170 304482 154226
rect 304538 154170 335078 154226
rect 335134 154170 335202 154226
rect 335258 154170 365798 154226
rect 365854 154170 365922 154226
rect 365978 154170 396518 154226
rect 396574 154170 396642 154226
rect 396698 154170 427238 154226
rect 427294 154170 427362 154226
rect 427418 154170 457958 154226
rect 458014 154170 458082 154226
rect 458138 154170 488678 154226
rect 488734 154170 488802 154226
rect 488858 154170 519398 154226
rect 519454 154170 519522 154226
rect 519578 154170 550118 154226
rect 550174 154170 550242 154226
rect 550298 154170 592914 154226
rect 592970 154170 593038 154226
rect 593094 154170 593162 154226
rect 593218 154170 593286 154226
rect 593342 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect -1916 154102 597980 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 27878 154102
rect 27934 154046 28002 154102
rect 28058 154046 58598 154102
rect 58654 154046 58722 154102
rect 58778 154046 89318 154102
rect 89374 154046 89442 154102
rect 89498 154046 120038 154102
rect 120094 154046 120162 154102
rect 120218 154046 150758 154102
rect 150814 154046 150882 154102
rect 150938 154046 181478 154102
rect 181534 154046 181602 154102
rect 181658 154046 212198 154102
rect 212254 154046 212322 154102
rect 212378 154046 242918 154102
rect 242974 154046 243042 154102
rect 243098 154046 273638 154102
rect 273694 154046 273762 154102
rect 273818 154046 304358 154102
rect 304414 154046 304482 154102
rect 304538 154046 335078 154102
rect 335134 154046 335202 154102
rect 335258 154046 365798 154102
rect 365854 154046 365922 154102
rect 365978 154046 396518 154102
rect 396574 154046 396642 154102
rect 396698 154046 427238 154102
rect 427294 154046 427362 154102
rect 427418 154046 457958 154102
rect 458014 154046 458082 154102
rect 458138 154046 488678 154102
rect 488734 154046 488802 154102
rect 488858 154046 519398 154102
rect 519454 154046 519522 154102
rect 519578 154046 550118 154102
rect 550174 154046 550242 154102
rect 550298 154046 592914 154102
rect 592970 154046 593038 154102
rect 593094 154046 593162 154102
rect 593218 154046 593286 154102
rect 593342 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect -1916 153978 597980 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 27878 153978
rect 27934 153922 28002 153978
rect 28058 153922 58598 153978
rect 58654 153922 58722 153978
rect 58778 153922 89318 153978
rect 89374 153922 89442 153978
rect 89498 153922 120038 153978
rect 120094 153922 120162 153978
rect 120218 153922 150758 153978
rect 150814 153922 150882 153978
rect 150938 153922 181478 153978
rect 181534 153922 181602 153978
rect 181658 153922 212198 153978
rect 212254 153922 212322 153978
rect 212378 153922 242918 153978
rect 242974 153922 243042 153978
rect 243098 153922 273638 153978
rect 273694 153922 273762 153978
rect 273818 153922 304358 153978
rect 304414 153922 304482 153978
rect 304538 153922 335078 153978
rect 335134 153922 335202 153978
rect 335258 153922 365798 153978
rect 365854 153922 365922 153978
rect 365978 153922 396518 153978
rect 396574 153922 396642 153978
rect 396698 153922 427238 153978
rect 427294 153922 427362 153978
rect 427418 153922 457958 153978
rect 458014 153922 458082 153978
rect 458138 153922 488678 153978
rect 488734 153922 488802 153978
rect 488858 153922 519398 153978
rect 519454 153922 519522 153978
rect 519578 153922 550118 153978
rect 550174 153922 550242 153978
rect 550298 153922 592914 153978
rect 592970 153922 593038 153978
rect 593094 153922 593162 153978
rect 593218 153922 593286 153978
rect 593342 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect -1916 153826 597980 153922
rect -1916 148350 597980 148446
rect -1916 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 5514 148350
rect 5570 148294 5638 148350
rect 5694 148294 5762 148350
rect 5818 148294 5886 148350
rect 5942 148294 12518 148350
rect 12574 148294 12642 148350
rect 12698 148294 43238 148350
rect 43294 148294 43362 148350
rect 43418 148294 73958 148350
rect 74014 148294 74082 148350
rect 74138 148294 104678 148350
rect 104734 148294 104802 148350
rect 104858 148294 135398 148350
rect 135454 148294 135522 148350
rect 135578 148294 166118 148350
rect 166174 148294 166242 148350
rect 166298 148294 196838 148350
rect 196894 148294 196962 148350
rect 197018 148294 227558 148350
rect 227614 148294 227682 148350
rect 227738 148294 258278 148350
rect 258334 148294 258402 148350
rect 258458 148294 288998 148350
rect 289054 148294 289122 148350
rect 289178 148294 319718 148350
rect 319774 148294 319842 148350
rect 319898 148294 350438 148350
rect 350494 148294 350562 148350
rect 350618 148294 381158 148350
rect 381214 148294 381282 148350
rect 381338 148294 411878 148350
rect 411934 148294 412002 148350
rect 412058 148294 442598 148350
rect 442654 148294 442722 148350
rect 442778 148294 473318 148350
rect 473374 148294 473442 148350
rect 473498 148294 504038 148350
rect 504094 148294 504162 148350
rect 504218 148294 534758 148350
rect 534814 148294 534882 148350
rect 534938 148294 565478 148350
rect 565534 148294 565602 148350
rect 565658 148294 589194 148350
rect 589250 148294 589318 148350
rect 589374 148294 589442 148350
rect 589498 148294 589566 148350
rect 589622 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597980 148350
rect -1916 148226 597980 148294
rect -1916 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 5514 148226
rect 5570 148170 5638 148226
rect 5694 148170 5762 148226
rect 5818 148170 5886 148226
rect 5942 148170 12518 148226
rect 12574 148170 12642 148226
rect 12698 148170 43238 148226
rect 43294 148170 43362 148226
rect 43418 148170 73958 148226
rect 74014 148170 74082 148226
rect 74138 148170 104678 148226
rect 104734 148170 104802 148226
rect 104858 148170 135398 148226
rect 135454 148170 135522 148226
rect 135578 148170 166118 148226
rect 166174 148170 166242 148226
rect 166298 148170 196838 148226
rect 196894 148170 196962 148226
rect 197018 148170 227558 148226
rect 227614 148170 227682 148226
rect 227738 148170 258278 148226
rect 258334 148170 258402 148226
rect 258458 148170 288998 148226
rect 289054 148170 289122 148226
rect 289178 148170 319718 148226
rect 319774 148170 319842 148226
rect 319898 148170 350438 148226
rect 350494 148170 350562 148226
rect 350618 148170 381158 148226
rect 381214 148170 381282 148226
rect 381338 148170 411878 148226
rect 411934 148170 412002 148226
rect 412058 148170 442598 148226
rect 442654 148170 442722 148226
rect 442778 148170 473318 148226
rect 473374 148170 473442 148226
rect 473498 148170 504038 148226
rect 504094 148170 504162 148226
rect 504218 148170 534758 148226
rect 534814 148170 534882 148226
rect 534938 148170 565478 148226
rect 565534 148170 565602 148226
rect 565658 148170 589194 148226
rect 589250 148170 589318 148226
rect 589374 148170 589442 148226
rect 589498 148170 589566 148226
rect 589622 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597980 148226
rect -1916 148102 597980 148170
rect -1916 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 5514 148102
rect 5570 148046 5638 148102
rect 5694 148046 5762 148102
rect 5818 148046 5886 148102
rect 5942 148046 12518 148102
rect 12574 148046 12642 148102
rect 12698 148046 43238 148102
rect 43294 148046 43362 148102
rect 43418 148046 73958 148102
rect 74014 148046 74082 148102
rect 74138 148046 104678 148102
rect 104734 148046 104802 148102
rect 104858 148046 135398 148102
rect 135454 148046 135522 148102
rect 135578 148046 166118 148102
rect 166174 148046 166242 148102
rect 166298 148046 196838 148102
rect 196894 148046 196962 148102
rect 197018 148046 227558 148102
rect 227614 148046 227682 148102
rect 227738 148046 258278 148102
rect 258334 148046 258402 148102
rect 258458 148046 288998 148102
rect 289054 148046 289122 148102
rect 289178 148046 319718 148102
rect 319774 148046 319842 148102
rect 319898 148046 350438 148102
rect 350494 148046 350562 148102
rect 350618 148046 381158 148102
rect 381214 148046 381282 148102
rect 381338 148046 411878 148102
rect 411934 148046 412002 148102
rect 412058 148046 442598 148102
rect 442654 148046 442722 148102
rect 442778 148046 473318 148102
rect 473374 148046 473442 148102
rect 473498 148046 504038 148102
rect 504094 148046 504162 148102
rect 504218 148046 534758 148102
rect 534814 148046 534882 148102
rect 534938 148046 565478 148102
rect 565534 148046 565602 148102
rect 565658 148046 589194 148102
rect 589250 148046 589318 148102
rect 589374 148046 589442 148102
rect 589498 148046 589566 148102
rect 589622 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597980 148102
rect -1916 147978 597980 148046
rect -1916 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 5514 147978
rect 5570 147922 5638 147978
rect 5694 147922 5762 147978
rect 5818 147922 5886 147978
rect 5942 147922 12518 147978
rect 12574 147922 12642 147978
rect 12698 147922 43238 147978
rect 43294 147922 43362 147978
rect 43418 147922 73958 147978
rect 74014 147922 74082 147978
rect 74138 147922 104678 147978
rect 104734 147922 104802 147978
rect 104858 147922 135398 147978
rect 135454 147922 135522 147978
rect 135578 147922 166118 147978
rect 166174 147922 166242 147978
rect 166298 147922 196838 147978
rect 196894 147922 196962 147978
rect 197018 147922 227558 147978
rect 227614 147922 227682 147978
rect 227738 147922 258278 147978
rect 258334 147922 258402 147978
rect 258458 147922 288998 147978
rect 289054 147922 289122 147978
rect 289178 147922 319718 147978
rect 319774 147922 319842 147978
rect 319898 147922 350438 147978
rect 350494 147922 350562 147978
rect 350618 147922 381158 147978
rect 381214 147922 381282 147978
rect 381338 147922 411878 147978
rect 411934 147922 412002 147978
rect 412058 147922 442598 147978
rect 442654 147922 442722 147978
rect 442778 147922 473318 147978
rect 473374 147922 473442 147978
rect 473498 147922 504038 147978
rect 504094 147922 504162 147978
rect 504218 147922 534758 147978
rect 534814 147922 534882 147978
rect 534938 147922 565478 147978
rect 565534 147922 565602 147978
rect 565658 147922 589194 147978
rect 589250 147922 589318 147978
rect 589374 147922 589442 147978
rect 589498 147922 589566 147978
rect 589622 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597980 147978
rect -1916 147826 597980 147922
rect -1916 136350 597980 136446
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 27878 136350
rect 27934 136294 28002 136350
rect 28058 136294 58598 136350
rect 58654 136294 58722 136350
rect 58778 136294 89318 136350
rect 89374 136294 89442 136350
rect 89498 136294 120038 136350
rect 120094 136294 120162 136350
rect 120218 136294 150758 136350
rect 150814 136294 150882 136350
rect 150938 136294 181478 136350
rect 181534 136294 181602 136350
rect 181658 136294 212198 136350
rect 212254 136294 212322 136350
rect 212378 136294 242918 136350
rect 242974 136294 243042 136350
rect 243098 136294 273638 136350
rect 273694 136294 273762 136350
rect 273818 136294 304358 136350
rect 304414 136294 304482 136350
rect 304538 136294 335078 136350
rect 335134 136294 335202 136350
rect 335258 136294 365798 136350
rect 365854 136294 365922 136350
rect 365978 136294 396518 136350
rect 396574 136294 396642 136350
rect 396698 136294 427238 136350
rect 427294 136294 427362 136350
rect 427418 136294 457958 136350
rect 458014 136294 458082 136350
rect 458138 136294 488678 136350
rect 488734 136294 488802 136350
rect 488858 136294 519398 136350
rect 519454 136294 519522 136350
rect 519578 136294 550118 136350
rect 550174 136294 550242 136350
rect 550298 136294 592914 136350
rect 592970 136294 593038 136350
rect 593094 136294 593162 136350
rect 593218 136294 593286 136350
rect 593342 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect -1916 136226 597980 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 27878 136226
rect 27934 136170 28002 136226
rect 28058 136170 58598 136226
rect 58654 136170 58722 136226
rect 58778 136170 89318 136226
rect 89374 136170 89442 136226
rect 89498 136170 120038 136226
rect 120094 136170 120162 136226
rect 120218 136170 150758 136226
rect 150814 136170 150882 136226
rect 150938 136170 181478 136226
rect 181534 136170 181602 136226
rect 181658 136170 212198 136226
rect 212254 136170 212322 136226
rect 212378 136170 242918 136226
rect 242974 136170 243042 136226
rect 243098 136170 273638 136226
rect 273694 136170 273762 136226
rect 273818 136170 304358 136226
rect 304414 136170 304482 136226
rect 304538 136170 335078 136226
rect 335134 136170 335202 136226
rect 335258 136170 365798 136226
rect 365854 136170 365922 136226
rect 365978 136170 396518 136226
rect 396574 136170 396642 136226
rect 396698 136170 427238 136226
rect 427294 136170 427362 136226
rect 427418 136170 457958 136226
rect 458014 136170 458082 136226
rect 458138 136170 488678 136226
rect 488734 136170 488802 136226
rect 488858 136170 519398 136226
rect 519454 136170 519522 136226
rect 519578 136170 550118 136226
rect 550174 136170 550242 136226
rect 550298 136170 592914 136226
rect 592970 136170 593038 136226
rect 593094 136170 593162 136226
rect 593218 136170 593286 136226
rect 593342 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect -1916 136102 597980 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 27878 136102
rect 27934 136046 28002 136102
rect 28058 136046 58598 136102
rect 58654 136046 58722 136102
rect 58778 136046 89318 136102
rect 89374 136046 89442 136102
rect 89498 136046 120038 136102
rect 120094 136046 120162 136102
rect 120218 136046 150758 136102
rect 150814 136046 150882 136102
rect 150938 136046 181478 136102
rect 181534 136046 181602 136102
rect 181658 136046 212198 136102
rect 212254 136046 212322 136102
rect 212378 136046 242918 136102
rect 242974 136046 243042 136102
rect 243098 136046 273638 136102
rect 273694 136046 273762 136102
rect 273818 136046 304358 136102
rect 304414 136046 304482 136102
rect 304538 136046 335078 136102
rect 335134 136046 335202 136102
rect 335258 136046 365798 136102
rect 365854 136046 365922 136102
rect 365978 136046 396518 136102
rect 396574 136046 396642 136102
rect 396698 136046 427238 136102
rect 427294 136046 427362 136102
rect 427418 136046 457958 136102
rect 458014 136046 458082 136102
rect 458138 136046 488678 136102
rect 488734 136046 488802 136102
rect 488858 136046 519398 136102
rect 519454 136046 519522 136102
rect 519578 136046 550118 136102
rect 550174 136046 550242 136102
rect 550298 136046 592914 136102
rect 592970 136046 593038 136102
rect 593094 136046 593162 136102
rect 593218 136046 593286 136102
rect 593342 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect -1916 135978 597980 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 27878 135978
rect 27934 135922 28002 135978
rect 28058 135922 58598 135978
rect 58654 135922 58722 135978
rect 58778 135922 89318 135978
rect 89374 135922 89442 135978
rect 89498 135922 120038 135978
rect 120094 135922 120162 135978
rect 120218 135922 150758 135978
rect 150814 135922 150882 135978
rect 150938 135922 181478 135978
rect 181534 135922 181602 135978
rect 181658 135922 212198 135978
rect 212254 135922 212322 135978
rect 212378 135922 242918 135978
rect 242974 135922 243042 135978
rect 243098 135922 273638 135978
rect 273694 135922 273762 135978
rect 273818 135922 304358 135978
rect 304414 135922 304482 135978
rect 304538 135922 335078 135978
rect 335134 135922 335202 135978
rect 335258 135922 365798 135978
rect 365854 135922 365922 135978
rect 365978 135922 396518 135978
rect 396574 135922 396642 135978
rect 396698 135922 427238 135978
rect 427294 135922 427362 135978
rect 427418 135922 457958 135978
rect 458014 135922 458082 135978
rect 458138 135922 488678 135978
rect 488734 135922 488802 135978
rect 488858 135922 519398 135978
rect 519454 135922 519522 135978
rect 519578 135922 550118 135978
rect 550174 135922 550242 135978
rect 550298 135922 592914 135978
rect 592970 135922 593038 135978
rect 593094 135922 593162 135978
rect 593218 135922 593286 135978
rect 593342 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect -1916 135826 597980 135922
rect -1916 130350 597980 130446
rect -1916 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 5514 130350
rect 5570 130294 5638 130350
rect 5694 130294 5762 130350
rect 5818 130294 5886 130350
rect 5942 130294 12518 130350
rect 12574 130294 12642 130350
rect 12698 130294 43238 130350
rect 43294 130294 43362 130350
rect 43418 130294 73958 130350
rect 74014 130294 74082 130350
rect 74138 130294 104678 130350
rect 104734 130294 104802 130350
rect 104858 130294 135398 130350
rect 135454 130294 135522 130350
rect 135578 130294 166118 130350
rect 166174 130294 166242 130350
rect 166298 130294 196838 130350
rect 196894 130294 196962 130350
rect 197018 130294 227558 130350
rect 227614 130294 227682 130350
rect 227738 130294 258278 130350
rect 258334 130294 258402 130350
rect 258458 130294 288998 130350
rect 289054 130294 289122 130350
rect 289178 130294 319718 130350
rect 319774 130294 319842 130350
rect 319898 130294 350438 130350
rect 350494 130294 350562 130350
rect 350618 130294 381158 130350
rect 381214 130294 381282 130350
rect 381338 130294 411878 130350
rect 411934 130294 412002 130350
rect 412058 130294 442598 130350
rect 442654 130294 442722 130350
rect 442778 130294 473318 130350
rect 473374 130294 473442 130350
rect 473498 130294 504038 130350
rect 504094 130294 504162 130350
rect 504218 130294 534758 130350
rect 534814 130294 534882 130350
rect 534938 130294 565478 130350
rect 565534 130294 565602 130350
rect 565658 130294 589194 130350
rect 589250 130294 589318 130350
rect 589374 130294 589442 130350
rect 589498 130294 589566 130350
rect 589622 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597980 130350
rect -1916 130226 597980 130294
rect -1916 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 5514 130226
rect 5570 130170 5638 130226
rect 5694 130170 5762 130226
rect 5818 130170 5886 130226
rect 5942 130170 12518 130226
rect 12574 130170 12642 130226
rect 12698 130170 43238 130226
rect 43294 130170 43362 130226
rect 43418 130170 73958 130226
rect 74014 130170 74082 130226
rect 74138 130170 104678 130226
rect 104734 130170 104802 130226
rect 104858 130170 135398 130226
rect 135454 130170 135522 130226
rect 135578 130170 166118 130226
rect 166174 130170 166242 130226
rect 166298 130170 196838 130226
rect 196894 130170 196962 130226
rect 197018 130170 227558 130226
rect 227614 130170 227682 130226
rect 227738 130170 258278 130226
rect 258334 130170 258402 130226
rect 258458 130170 288998 130226
rect 289054 130170 289122 130226
rect 289178 130170 319718 130226
rect 319774 130170 319842 130226
rect 319898 130170 350438 130226
rect 350494 130170 350562 130226
rect 350618 130170 381158 130226
rect 381214 130170 381282 130226
rect 381338 130170 411878 130226
rect 411934 130170 412002 130226
rect 412058 130170 442598 130226
rect 442654 130170 442722 130226
rect 442778 130170 473318 130226
rect 473374 130170 473442 130226
rect 473498 130170 504038 130226
rect 504094 130170 504162 130226
rect 504218 130170 534758 130226
rect 534814 130170 534882 130226
rect 534938 130170 565478 130226
rect 565534 130170 565602 130226
rect 565658 130170 589194 130226
rect 589250 130170 589318 130226
rect 589374 130170 589442 130226
rect 589498 130170 589566 130226
rect 589622 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597980 130226
rect -1916 130102 597980 130170
rect -1916 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 5514 130102
rect 5570 130046 5638 130102
rect 5694 130046 5762 130102
rect 5818 130046 5886 130102
rect 5942 130046 12518 130102
rect 12574 130046 12642 130102
rect 12698 130046 43238 130102
rect 43294 130046 43362 130102
rect 43418 130046 73958 130102
rect 74014 130046 74082 130102
rect 74138 130046 104678 130102
rect 104734 130046 104802 130102
rect 104858 130046 135398 130102
rect 135454 130046 135522 130102
rect 135578 130046 166118 130102
rect 166174 130046 166242 130102
rect 166298 130046 196838 130102
rect 196894 130046 196962 130102
rect 197018 130046 227558 130102
rect 227614 130046 227682 130102
rect 227738 130046 258278 130102
rect 258334 130046 258402 130102
rect 258458 130046 288998 130102
rect 289054 130046 289122 130102
rect 289178 130046 319718 130102
rect 319774 130046 319842 130102
rect 319898 130046 350438 130102
rect 350494 130046 350562 130102
rect 350618 130046 381158 130102
rect 381214 130046 381282 130102
rect 381338 130046 411878 130102
rect 411934 130046 412002 130102
rect 412058 130046 442598 130102
rect 442654 130046 442722 130102
rect 442778 130046 473318 130102
rect 473374 130046 473442 130102
rect 473498 130046 504038 130102
rect 504094 130046 504162 130102
rect 504218 130046 534758 130102
rect 534814 130046 534882 130102
rect 534938 130046 565478 130102
rect 565534 130046 565602 130102
rect 565658 130046 589194 130102
rect 589250 130046 589318 130102
rect 589374 130046 589442 130102
rect 589498 130046 589566 130102
rect 589622 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597980 130102
rect -1916 129978 597980 130046
rect -1916 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 5514 129978
rect 5570 129922 5638 129978
rect 5694 129922 5762 129978
rect 5818 129922 5886 129978
rect 5942 129922 12518 129978
rect 12574 129922 12642 129978
rect 12698 129922 43238 129978
rect 43294 129922 43362 129978
rect 43418 129922 73958 129978
rect 74014 129922 74082 129978
rect 74138 129922 104678 129978
rect 104734 129922 104802 129978
rect 104858 129922 135398 129978
rect 135454 129922 135522 129978
rect 135578 129922 166118 129978
rect 166174 129922 166242 129978
rect 166298 129922 196838 129978
rect 196894 129922 196962 129978
rect 197018 129922 227558 129978
rect 227614 129922 227682 129978
rect 227738 129922 258278 129978
rect 258334 129922 258402 129978
rect 258458 129922 288998 129978
rect 289054 129922 289122 129978
rect 289178 129922 319718 129978
rect 319774 129922 319842 129978
rect 319898 129922 350438 129978
rect 350494 129922 350562 129978
rect 350618 129922 381158 129978
rect 381214 129922 381282 129978
rect 381338 129922 411878 129978
rect 411934 129922 412002 129978
rect 412058 129922 442598 129978
rect 442654 129922 442722 129978
rect 442778 129922 473318 129978
rect 473374 129922 473442 129978
rect 473498 129922 504038 129978
rect 504094 129922 504162 129978
rect 504218 129922 534758 129978
rect 534814 129922 534882 129978
rect 534938 129922 565478 129978
rect 565534 129922 565602 129978
rect 565658 129922 589194 129978
rect 589250 129922 589318 129978
rect 589374 129922 589442 129978
rect 589498 129922 589566 129978
rect 589622 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597980 129978
rect -1916 129826 597980 129922
rect -1916 118350 597980 118446
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 27878 118350
rect 27934 118294 28002 118350
rect 28058 118294 58598 118350
rect 58654 118294 58722 118350
rect 58778 118294 89318 118350
rect 89374 118294 89442 118350
rect 89498 118294 120038 118350
rect 120094 118294 120162 118350
rect 120218 118294 150758 118350
rect 150814 118294 150882 118350
rect 150938 118294 181478 118350
rect 181534 118294 181602 118350
rect 181658 118294 212198 118350
rect 212254 118294 212322 118350
rect 212378 118294 242918 118350
rect 242974 118294 243042 118350
rect 243098 118294 273638 118350
rect 273694 118294 273762 118350
rect 273818 118294 304358 118350
rect 304414 118294 304482 118350
rect 304538 118294 335078 118350
rect 335134 118294 335202 118350
rect 335258 118294 365798 118350
rect 365854 118294 365922 118350
rect 365978 118294 396518 118350
rect 396574 118294 396642 118350
rect 396698 118294 427238 118350
rect 427294 118294 427362 118350
rect 427418 118294 457958 118350
rect 458014 118294 458082 118350
rect 458138 118294 488678 118350
rect 488734 118294 488802 118350
rect 488858 118294 519398 118350
rect 519454 118294 519522 118350
rect 519578 118294 550118 118350
rect 550174 118294 550242 118350
rect 550298 118294 592914 118350
rect 592970 118294 593038 118350
rect 593094 118294 593162 118350
rect 593218 118294 593286 118350
rect 593342 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect -1916 118226 597980 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 27878 118226
rect 27934 118170 28002 118226
rect 28058 118170 58598 118226
rect 58654 118170 58722 118226
rect 58778 118170 89318 118226
rect 89374 118170 89442 118226
rect 89498 118170 120038 118226
rect 120094 118170 120162 118226
rect 120218 118170 150758 118226
rect 150814 118170 150882 118226
rect 150938 118170 181478 118226
rect 181534 118170 181602 118226
rect 181658 118170 212198 118226
rect 212254 118170 212322 118226
rect 212378 118170 242918 118226
rect 242974 118170 243042 118226
rect 243098 118170 273638 118226
rect 273694 118170 273762 118226
rect 273818 118170 304358 118226
rect 304414 118170 304482 118226
rect 304538 118170 335078 118226
rect 335134 118170 335202 118226
rect 335258 118170 365798 118226
rect 365854 118170 365922 118226
rect 365978 118170 396518 118226
rect 396574 118170 396642 118226
rect 396698 118170 427238 118226
rect 427294 118170 427362 118226
rect 427418 118170 457958 118226
rect 458014 118170 458082 118226
rect 458138 118170 488678 118226
rect 488734 118170 488802 118226
rect 488858 118170 519398 118226
rect 519454 118170 519522 118226
rect 519578 118170 550118 118226
rect 550174 118170 550242 118226
rect 550298 118170 592914 118226
rect 592970 118170 593038 118226
rect 593094 118170 593162 118226
rect 593218 118170 593286 118226
rect 593342 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect -1916 118102 597980 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 27878 118102
rect 27934 118046 28002 118102
rect 28058 118046 58598 118102
rect 58654 118046 58722 118102
rect 58778 118046 89318 118102
rect 89374 118046 89442 118102
rect 89498 118046 120038 118102
rect 120094 118046 120162 118102
rect 120218 118046 150758 118102
rect 150814 118046 150882 118102
rect 150938 118046 181478 118102
rect 181534 118046 181602 118102
rect 181658 118046 212198 118102
rect 212254 118046 212322 118102
rect 212378 118046 242918 118102
rect 242974 118046 243042 118102
rect 243098 118046 273638 118102
rect 273694 118046 273762 118102
rect 273818 118046 304358 118102
rect 304414 118046 304482 118102
rect 304538 118046 335078 118102
rect 335134 118046 335202 118102
rect 335258 118046 365798 118102
rect 365854 118046 365922 118102
rect 365978 118046 396518 118102
rect 396574 118046 396642 118102
rect 396698 118046 427238 118102
rect 427294 118046 427362 118102
rect 427418 118046 457958 118102
rect 458014 118046 458082 118102
rect 458138 118046 488678 118102
rect 488734 118046 488802 118102
rect 488858 118046 519398 118102
rect 519454 118046 519522 118102
rect 519578 118046 550118 118102
rect 550174 118046 550242 118102
rect 550298 118046 592914 118102
rect 592970 118046 593038 118102
rect 593094 118046 593162 118102
rect 593218 118046 593286 118102
rect 593342 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect -1916 117978 597980 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 27878 117978
rect 27934 117922 28002 117978
rect 28058 117922 58598 117978
rect 58654 117922 58722 117978
rect 58778 117922 89318 117978
rect 89374 117922 89442 117978
rect 89498 117922 120038 117978
rect 120094 117922 120162 117978
rect 120218 117922 150758 117978
rect 150814 117922 150882 117978
rect 150938 117922 181478 117978
rect 181534 117922 181602 117978
rect 181658 117922 212198 117978
rect 212254 117922 212322 117978
rect 212378 117922 242918 117978
rect 242974 117922 243042 117978
rect 243098 117922 273638 117978
rect 273694 117922 273762 117978
rect 273818 117922 304358 117978
rect 304414 117922 304482 117978
rect 304538 117922 335078 117978
rect 335134 117922 335202 117978
rect 335258 117922 365798 117978
rect 365854 117922 365922 117978
rect 365978 117922 396518 117978
rect 396574 117922 396642 117978
rect 396698 117922 427238 117978
rect 427294 117922 427362 117978
rect 427418 117922 457958 117978
rect 458014 117922 458082 117978
rect 458138 117922 488678 117978
rect 488734 117922 488802 117978
rect 488858 117922 519398 117978
rect 519454 117922 519522 117978
rect 519578 117922 550118 117978
rect 550174 117922 550242 117978
rect 550298 117922 592914 117978
rect 592970 117922 593038 117978
rect 593094 117922 593162 117978
rect 593218 117922 593286 117978
rect 593342 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect -1916 117826 597980 117922
rect -1916 112350 597980 112446
rect -1916 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 5514 112350
rect 5570 112294 5638 112350
rect 5694 112294 5762 112350
rect 5818 112294 5886 112350
rect 5942 112294 12518 112350
rect 12574 112294 12642 112350
rect 12698 112294 43238 112350
rect 43294 112294 43362 112350
rect 43418 112294 73958 112350
rect 74014 112294 74082 112350
rect 74138 112294 104678 112350
rect 104734 112294 104802 112350
rect 104858 112294 135398 112350
rect 135454 112294 135522 112350
rect 135578 112294 166118 112350
rect 166174 112294 166242 112350
rect 166298 112294 196838 112350
rect 196894 112294 196962 112350
rect 197018 112294 227558 112350
rect 227614 112294 227682 112350
rect 227738 112294 258278 112350
rect 258334 112294 258402 112350
rect 258458 112294 288998 112350
rect 289054 112294 289122 112350
rect 289178 112294 319718 112350
rect 319774 112294 319842 112350
rect 319898 112294 350438 112350
rect 350494 112294 350562 112350
rect 350618 112294 381158 112350
rect 381214 112294 381282 112350
rect 381338 112294 411878 112350
rect 411934 112294 412002 112350
rect 412058 112294 442598 112350
rect 442654 112294 442722 112350
rect 442778 112294 473318 112350
rect 473374 112294 473442 112350
rect 473498 112294 504038 112350
rect 504094 112294 504162 112350
rect 504218 112294 534758 112350
rect 534814 112294 534882 112350
rect 534938 112294 565478 112350
rect 565534 112294 565602 112350
rect 565658 112294 589194 112350
rect 589250 112294 589318 112350
rect 589374 112294 589442 112350
rect 589498 112294 589566 112350
rect 589622 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597980 112350
rect -1916 112226 597980 112294
rect -1916 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 5514 112226
rect 5570 112170 5638 112226
rect 5694 112170 5762 112226
rect 5818 112170 5886 112226
rect 5942 112170 12518 112226
rect 12574 112170 12642 112226
rect 12698 112170 43238 112226
rect 43294 112170 43362 112226
rect 43418 112170 73958 112226
rect 74014 112170 74082 112226
rect 74138 112170 104678 112226
rect 104734 112170 104802 112226
rect 104858 112170 135398 112226
rect 135454 112170 135522 112226
rect 135578 112170 166118 112226
rect 166174 112170 166242 112226
rect 166298 112170 196838 112226
rect 196894 112170 196962 112226
rect 197018 112170 227558 112226
rect 227614 112170 227682 112226
rect 227738 112170 258278 112226
rect 258334 112170 258402 112226
rect 258458 112170 288998 112226
rect 289054 112170 289122 112226
rect 289178 112170 319718 112226
rect 319774 112170 319842 112226
rect 319898 112170 350438 112226
rect 350494 112170 350562 112226
rect 350618 112170 381158 112226
rect 381214 112170 381282 112226
rect 381338 112170 411878 112226
rect 411934 112170 412002 112226
rect 412058 112170 442598 112226
rect 442654 112170 442722 112226
rect 442778 112170 473318 112226
rect 473374 112170 473442 112226
rect 473498 112170 504038 112226
rect 504094 112170 504162 112226
rect 504218 112170 534758 112226
rect 534814 112170 534882 112226
rect 534938 112170 565478 112226
rect 565534 112170 565602 112226
rect 565658 112170 589194 112226
rect 589250 112170 589318 112226
rect 589374 112170 589442 112226
rect 589498 112170 589566 112226
rect 589622 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597980 112226
rect -1916 112102 597980 112170
rect -1916 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 5514 112102
rect 5570 112046 5638 112102
rect 5694 112046 5762 112102
rect 5818 112046 5886 112102
rect 5942 112046 12518 112102
rect 12574 112046 12642 112102
rect 12698 112046 43238 112102
rect 43294 112046 43362 112102
rect 43418 112046 73958 112102
rect 74014 112046 74082 112102
rect 74138 112046 104678 112102
rect 104734 112046 104802 112102
rect 104858 112046 135398 112102
rect 135454 112046 135522 112102
rect 135578 112046 166118 112102
rect 166174 112046 166242 112102
rect 166298 112046 196838 112102
rect 196894 112046 196962 112102
rect 197018 112046 227558 112102
rect 227614 112046 227682 112102
rect 227738 112046 258278 112102
rect 258334 112046 258402 112102
rect 258458 112046 288998 112102
rect 289054 112046 289122 112102
rect 289178 112046 319718 112102
rect 319774 112046 319842 112102
rect 319898 112046 350438 112102
rect 350494 112046 350562 112102
rect 350618 112046 381158 112102
rect 381214 112046 381282 112102
rect 381338 112046 411878 112102
rect 411934 112046 412002 112102
rect 412058 112046 442598 112102
rect 442654 112046 442722 112102
rect 442778 112046 473318 112102
rect 473374 112046 473442 112102
rect 473498 112046 504038 112102
rect 504094 112046 504162 112102
rect 504218 112046 534758 112102
rect 534814 112046 534882 112102
rect 534938 112046 565478 112102
rect 565534 112046 565602 112102
rect 565658 112046 589194 112102
rect 589250 112046 589318 112102
rect 589374 112046 589442 112102
rect 589498 112046 589566 112102
rect 589622 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597980 112102
rect -1916 111978 597980 112046
rect -1916 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 5514 111978
rect 5570 111922 5638 111978
rect 5694 111922 5762 111978
rect 5818 111922 5886 111978
rect 5942 111922 12518 111978
rect 12574 111922 12642 111978
rect 12698 111922 43238 111978
rect 43294 111922 43362 111978
rect 43418 111922 73958 111978
rect 74014 111922 74082 111978
rect 74138 111922 104678 111978
rect 104734 111922 104802 111978
rect 104858 111922 135398 111978
rect 135454 111922 135522 111978
rect 135578 111922 166118 111978
rect 166174 111922 166242 111978
rect 166298 111922 196838 111978
rect 196894 111922 196962 111978
rect 197018 111922 227558 111978
rect 227614 111922 227682 111978
rect 227738 111922 258278 111978
rect 258334 111922 258402 111978
rect 258458 111922 288998 111978
rect 289054 111922 289122 111978
rect 289178 111922 319718 111978
rect 319774 111922 319842 111978
rect 319898 111922 350438 111978
rect 350494 111922 350562 111978
rect 350618 111922 381158 111978
rect 381214 111922 381282 111978
rect 381338 111922 411878 111978
rect 411934 111922 412002 111978
rect 412058 111922 442598 111978
rect 442654 111922 442722 111978
rect 442778 111922 473318 111978
rect 473374 111922 473442 111978
rect 473498 111922 504038 111978
rect 504094 111922 504162 111978
rect 504218 111922 534758 111978
rect 534814 111922 534882 111978
rect 534938 111922 565478 111978
rect 565534 111922 565602 111978
rect 565658 111922 589194 111978
rect 589250 111922 589318 111978
rect 589374 111922 589442 111978
rect 589498 111922 589566 111978
rect 589622 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597980 111978
rect -1916 111826 597980 111922
rect -1916 100350 597980 100446
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 27878 100350
rect 27934 100294 28002 100350
rect 28058 100294 58598 100350
rect 58654 100294 58722 100350
rect 58778 100294 89318 100350
rect 89374 100294 89442 100350
rect 89498 100294 120038 100350
rect 120094 100294 120162 100350
rect 120218 100294 150758 100350
rect 150814 100294 150882 100350
rect 150938 100294 181478 100350
rect 181534 100294 181602 100350
rect 181658 100294 212198 100350
rect 212254 100294 212322 100350
rect 212378 100294 242918 100350
rect 242974 100294 243042 100350
rect 243098 100294 273638 100350
rect 273694 100294 273762 100350
rect 273818 100294 304358 100350
rect 304414 100294 304482 100350
rect 304538 100294 335078 100350
rect 335134 100294 335202 100350
rect 335258 100294 365798 100350
rect 365854 100294 365922 100350
rect 365978 100294 396518 100350
rect 396574 100294 396642 100350
rect 396698 100294 427238 100350
rect 427294 100294 427362 100350
rect 427418 100294 457958 100350
rect 458014 100294 458082 100350
rect 458138 100294 488678 100350
rect 488734 100294 488802 100350
rect 488858 100294 519398 100350
rect 519454 100294 519522 100350
rect 519578 100294 550118 100350
rect 550174 100294 550242 100350
rect 550298 100294 592914 100350
rect 592970 100294 593038 100350
rect 593094 100294 593162 100350
rect 593218 100294 593286 100350
rect 593342 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect -1916 100226 597980 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 27878 100226
rect 27934 100170 28002 100226
rect 28058 100170 58598 100226
rect 58654 100170 58722 100226
rect 58778 100170 89318 100226
rect 89374 100170 89442 100226
rect 89498 100170 120038 100226
rect 120094 100170 120162 100226
rect 120218 100170 150758 100226
rect 150814 100170 150882 100226
rect 150938 100170 181478 100226
rect 181534 100170 181602 100226
rect 181658 100170 212198 100226
rect 212254 100170 212322 100226
rect 212378 100170 242918 100226
rect 242974 100170 243042 100226
rect 243098 100170 273638 100226
rect 273694 100170 273762 100226
rect 273818 100170 304358 100226
rect 304414 100170 304482 100226
rect 304538 100170 335078 100226
rect 335134 100170 335202 100226
rect 335258 100170 365798 100226
rect 365854 100170 365922 100226
rect 365978 100170 396518 100226
rect 396574 100170 396642 100226
rect 396698 100170 427238 100226
rect 427294 100170 427362 100226
rect 427418 100170 457958 100226
rect 458014 100170 458082 100226
rect 458138 100170 488678 100226
rect 488734 100170 488802 100226
rect 488858 100170 519398 100226
rect 519454 100170 519522 100226
rect 519578 100170 550118 100226
rect 550174 100170 550242 100226
rect 550298 100170 592914 100226
rect 592970 100170 593038 100226
rect 593094 100170 593162 100226
rect 593218 100170 593286 100226
rect 593342 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect -1916 100102 597980 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 27878 100102
rect 27934 100046 28002 100102
rect 28058 100046 58598 100102
rect 58654 100046 58722 100102
rect 58778 100046 89318 100102
rect 89374 100046 89442 100102
rect 89498 100046 120038 100102
rect 120094 100046 120162 100102
rect 120218 100046 150758 100102
rect 150814 100046 150882 100102
rect 150938 100046 181478 100102
rect 181534 100046 181602 100102
rect 181658 100046 212198 100102
rect 212254 100046 212322 100102
rect 212378 100046 242918 100102
rect 242974 100046 243042 100102
rect 243098 100046 273638 100102
rect 273694 100046 273762 100102
rect 273818 100046 304358 100102
rect 304414 100046 304482 100102
rect 304538 100046 335078 100102
rect 335134 100046 335202 100102
rect 335258 100046 365798 100102
rect 365854 100046 365922 100102
rect 365978 100046 396518 100102
rect 396574 100046 396642 100102
rect 396698 100046 427238 100102
rect 427294 100046 427362 100102
rect 427418 100046 457958 100102
rect 458014 100046 458082 100102
rect 458138 100046 488678 100102
rect 488734 100046 488802 100102
rect 488858 100046 519398 100102
rect 519454 100046 519522 100102
rect 519578 100046 550118 100102
rect 550174 100046 550242 100102
rect 550298 100046 592914 100102
rect 592970 100046 593038 100102
rect 593094 100046 593162 100102
rect 593218 100046 593286 100102
rect 593342 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect -1916 99978 597980 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 27878 99978
rect 27934 99922 28002 99978
rect 28058 99922 58598 99978
rect 58654 99922 58722 99978
rect 58778 99922 89318 99978
rect 89374 99922 89442 99978
rect 89498 99922 120038 99978
rect 120094 99922 120162 99978
rect 120218 99922 150758 99978
rect 150814 99922 150882 99978
rect 150938 99922 181478 99978
rect 181534 99922 181602 99978
rect 181658 99922 212198 99978
rect 212254 99922 212322 99978
rect 212378 99922 242918 99978
rect 242974 99922 243042 99978
rect 243098 99922 273638 99978
rect 273694 99922 273762 99978
rect 273818 99922 304358 99978
rect 304414 99922 304482 99978
rect 304538 99922 335078 99978
rect 335134 99922 335202 99978
rect 335258 99922 365798 99978
rect 365854 99922 365922 99978
rect 365978 99922 396518 99978
rect 396574 99922 396642 99978
rect 396698 99922 427238 99978
rect 427294 99922 427362 99978
rect 427418 99922 457958 99978
rect 458014 99922 458082 99978
rect 458138 99922 488678 99978
rect 488734 99922 488802 99978
rect 488858 99922 519398 99978
rect 519454 99922 519522 99978
rect 519578 99922 550118 99978
rect 550174 99922 550242 99978
rect 550298 99922 592914 99978
rect 592970 99922 593038 99978
rect 593094 99922 593162 99978
rect 593218 99922 593286 99978
rect 593342 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect -1916 99826 597980 99922
rect -1916 94350 597980 94446
rect -1916 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 5514 94350
rect 5570 94294 5638 94350
rect 5694 94294 5762 94350
rect 5818 94294 5886 94350
rect 5942 94294 12518 94350
rect 12574 94294 12642 94350
rect 12698 94294 43238 94350
rect 43294 94294 43362 94350
rect 43418 94294 73958 94350
rect 74014 94294 74082 94350
rect 74138 94294 104678 94350
rect 104734 94294 104802 94350
rect 104858 94294 135398 94350
rect 135454 94294 135522 94350
rect 135578 94294 166118 94350
rect 166174 94294 166242 94350
rect 166298 94294 196838 94350
rect 196894 94294 196962 94350
rect 197018 94294 227558 94350
rect 227614 94294 227682 94350
rect 227738 94294 258278 94350
rect 258334 94294 258402 94350
rect 258458 94294 288998 94350
rect 289054 94294 289122 94350
rect 289178 94294 319718 94350
rect 319774 94294 319842 94350
rect 319898 94294 350438 94350
rect 350494 94294 350562 94350
rect 350618 94294 381158 94350
rect 381214 94294 381282 94350
rect 381338 94294 411878 94350
rect 411934 94294 412002 94350
rect 412058 94294 442598 94350
rect 442654 94294 442722 94350
rect 442778 94294 473318 94350
rect 473374 94294 473442 94350
rect 473498 94294 504038 94350
rect 504094 94294 504162 94350
rect 504218 94294 534758 94350
rect 534814 94294 534882 94350
rect 534938 94294 565478 94350
rect 565534 94294 565602 94350
rect 565658 94294 589194 94350
rect 589250 94294 589318 94350
rect 589374 94294 589442 94350
rect 589498 94294 589566 94350
rect 589622 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597980 94350
rect -1916 94226 597980 94294
rect -1916 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 5514 94226
rect 5570 94170 5638 94226
rect 5694 94170 5762 94226
rect 5818 94170 5886 94226
rect 5942 94170 12518 94226
rect 12574 94170 12642 94226
rect 12698 94170 43238 94226
rect 43294 94170 43362 94226
rect 43418 94170 73958 94226
rect 74014 94170 74082 94226
rect 74138 94170 104678 94226
rect 104734 94170 104802 94226
rect 104858 94170 135398 94226
rect 135454 94170 135522 94226
rect 135578 94170 166118 94226
rect 166174 94170 166242 94226
rect 166298 94170 196838 94226
rect 196894 94170 196962 94226
rect 197018 94170 227558 94226
rect 227614 94170 227682 94226
rect 227738 94170 258278 94226
rect 258334 94170 258402 94226
rect 258458 94170 288998 94226
rect 289054 94170 289122 94226
rect 289178 94170 319718 94226
rect 319774 94170 319842 94226
rect 319898 94170 350438 94226
rect 350494 94170 350562 94226
rect 350618 94170 381158 94226
rect 381214 94170 381282 94226
rect 381338 94170 411878 94226
rect 411934 94170 412002 94226
rect 412058 94170 442598 94226
rect 442654 94170 442722 94226
rect 442778 94170 473318 94226
rect 473374 94170 473442 94226
rect 473498 94170 504038 94226
rect 504094 94170 504162 94226
rect 504218 94170 534758 94226
rect 534814 94170 534882 94226
rect 534938 94170 565478 94226
rect 565534 94170 565602 94226
rect 565658 94170 589194 94226
rect 589250 94170 589318 94226
rect 589374 94170 589442 94226
rect 589498 94170 589566 94226
rect 589622 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597980 94226
rect -1916 94102 597980 94170
rect -1916 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 5514 94102
rect 5570 94046 5638 94102
rect 5694 94046 5762 94102
rect 5818 94046 5886 94102
rect 5942 94046 12518 94102
rect 12574 94046 12642 94102
rect 12698 94046 43238 94102
rect 43294 94046 43362 94102
rect 43418 94046 73958 94102
rect 74014 94046 74082 94102
rect 74138 94046 104678 94102
rect 104734 94046 104802 94102
rect 104858 94046 135398 94102
rect 135454 94046 135522 94102
rect 135578 94046 166118 94102
rect 166174 94046 166242 94102
rect 166298 94046 196838 94102
rect 196894 94046 196962 94102
rect 197018 94046 227558 94102
rect 227614 94046 227682 94102
rect 227738 94046 258278 94102
rect 258334 94046 258402 94102
rect 258458 94046 288998 94102
rect 289054 94046 289122 94102
rect 289178 94046 319718 94102
rect 319774 94046 319842 94102
rect 319898 94046 350438 94102
rect 350494 94046 350562 94102
rect 350618 94046 381158 94102
rect 381214 94046 381282 94102
rect 381338 94046 411878 94102
rect 411934 94046 412002 94102
rect 412058 94046 442598 94102
rect 442654 94046 442722 94102
rect 442778 94046 473318 94102
rect 473374 94046 473442 94102
rect 473498 94046 504038 94102
rect 504094 94046 504162 94102
rect 504218 94046 534758 94102
rect 534814 94046 534882 94102
rect 534938 94046 565478 94102
rect 565534 94046 565602 94102
rect 565658 94046 589194 94102
rect 589250 94046 589318 94102
rect 589374 94046 589442 94102
rect 589498 94046 589566 94102
rect 589622 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597980 94102
rect -1916 93978 597980 94046
rect -1916 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 5514 93978
rect 5570 93922 5638 93978
rect 5694 93922 5762 93978
rect 5818 93922 5886 93978
rect 5942 93922 12518 93978
rect 12574 93922 12642 93978
rect 12698 93922 43238 93978
rect 43294 93922 43362 93978
rect 43418 93922 73958 93978
rect 74014 93922 74082 93978
rect 74138 93922 104678 93978
rect 104734 93922 104802 93978
rect 104858 93922 135398 93978
rect 135454 93922 135522 93978
rect 135578 93922 166118 93978
rect 166174 93922 166242 93978
rect 166298 93922 196838 93978
rect 196894 93922 196962 93978
rect 197018 93922 227558 93978
rect 227614 93922 227682 93978
rect 227738 93922 258278 93978
rect 258334 93922 258402 93978
rect 258458 93922 288998 93978
rect 289054 93922 289122 93978
rect 289178 93922 319718 93978
rect 319774 93922 319842 93978
rect 319898 93922 350438 93978
rect 350494 93922 350562 93978
rect 350618 93922 381158 93978
rect 381214 93922 381282 93978
rect 381338 93922 411878 93978
rect 411934 93922 412002 93978
rect 412058 93922 442598 93978
rect 442654 93922 442722 93978
rect 442778 93922 473318 93978
rect 473374 93922 473442 93978
rect 473498 93922 504038 93978
rect 504094 93922 504162 93978
rect 504218 93922 534758 93978
rect 534814 93922 534882 93978
rect 534938 93922 565478 93978
rect 565534 93922 565602 93978
rect 565658 93922 589194 93978
rect 589250 93922 589318 93978
rect 589374 93922 589442 93978
rect 589498 93922 589566 93978
rect 589622 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597980 93978
rect -1916 93826 597980 93922
rect -1916 82350 597980 82446
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 27878 82350
rect 27934 82294 28002 82350
rect 28058 82294 58598 82350
rect 58654 82294 58722 82350
rect 58778 82294 89318 82350
rect 89374 82294 89442 82350
rect 89498 82294 120038 82350
rect 120094 82294 120162 82350
rect 120218 82294 150758 82350
rect 150814 82294 150882 82350
rect 150938 82294 181478 82350
rect 181534 82294 181602 82350
rect 181658 82294 212198 82350
rect 212254 82294 212322 82350
rect 212378 82294 242918 82350
rect 242974 82294 243042 82350
rect 243098 82294 273638 82350
rect 273694 82294 273762 82350
rect 273818 82294 304358 82350
rect 304414 82294 304482 82350
rect 304538 82294 335078 82350
rect 335134 82294 335202 82350
rect 335258 82294 365798 82350
rect 365854 82294 365922 82350
rect 365978 82294 396518 82350
rect 396574 82294 396642 82350
rect 396698 82294 427238 82350
rect 427294 82294 427362 82350
rect 427418 82294 457958 82350
rect 458014 82294 458082 82350
rect 458138 82294 488678 82350
rect 488734 82294 488802 82350
rect 488858 82294 519398 82350
rect 519454 82294 519522 82350
rect 519578 82294 550118 82350
rect 550174 82294 550242 82350
rect 550298 82294 592914 82350
rect 592970 82294 593038 82350
rect 593094 82294 593162 82350
rect 593218 82294 593286 82350
rect 593342 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect -1916 82226 597980 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 27878 82226
rect 27934 82170 28002 82226
rect 28058 82170 58598 82226
rect 58654 82170 58722 82226
rect 58778 82170 89318 82226
rect 89374 82170 89442 82226
rect 89498 82170 120038 82226
rect 120094 82170 120162 82226
rect 120218 82170 150758 82226
rect 150814 82170 150882 82226
rect 150938 82170 181478 82226
rect 181534 82170 181602 82226
rect 181658 82170 212198 82226
rect 212254 82170 212322 82226
rect 212378 82170 242918 82226
rect 242974 82170 243042 82226
rect 243098 82170 273638 82226
rect 273694 82170 273762 82226
rect 273818 82170 304358 82226
rect 304414 82170 304482 82226
rect 304538 82170 335078 82226
rect 335134 82170 335202 82226
rect 335258 82170 365798 82226
rect 365854 82170 365922 82226
rect 365978 82170 396518 82226
rect 396574 82170 396642 82226
rect 396698 82170 427238 82226
rect 427294 82170 427362 82226
rect 427418 82170 457958 82226
rect 458014 82170 458082 82226
rect 458138 82170 488678 82226
rect 488734 82170 488802 82226
rect 488858 82170 519398 82226
rect 519454 82170 519522 82226
rect 519578 82170 550118 82226
rect 550174 82170 550242 82226
rect 550298 82170 592914 82226
rect 592970 82170 593038 82226
rect 593094 82170 593162 82226
rect 593218 82170 593286 82226
rect 593342 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect -1916 82102 597980 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 27878 82102
rect 27934 82046 28002 82102
rect 28058 82046 58598 82102
rect 58654 82046 58722 82102
rect 58778 82046 89318 82102
rect 89374 82046 89442 82102
rect 89498 82046 120038 82102
rect 120094 82046 120162 82102
rect 120218 82046 150758 82102
rect 150814 82046 150882 82102
rect 150938 82046 181478 82102
rect 181534 82046 181602 82102
rect 181658 82046 212198 82102
rect 212254 82046 212322 82102
rect 212378 82046 242918 82102
rect 242974 82046 243042 82102
rect 243098 82046 273638 82102
rect 273694 82046 273762 82102
rect 273818 82046 304358 82102
rect 304414 82046 304482 82102
rect 304538 82046 335078 82102
rect 335134 82046 335202 82102
rect 335258 82046 365798 82102
rect 365854 82046 365922 82102
rect 365978 82046 396518 82102
rect 396574 82046 396642 82102
rect 396698 82046 427238 82102
rect 427294 82046 427362 82102
rect 427418 82046 457958 82102
rect 458014 82046 458082 82102
rect 458138 82046 488678 82102
rect 488734 82046 488802 82102
rect 488858 82046 519398 82102
rect 519454 82046 519522 82102
rect 519578 82046 550118 82102
rect 550174 82046 550242 82102
rect 550298 82046 592914 82102
rect 592970 82046 593038 82102
rect 593094 82046 593162 82102
rect 593218 82046 593286 82102
rect 593342 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect -1916 81978 597980 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 27878 81978
rect 27934 81922 28002 81978
rect 28058 81922 58598 81978
rect 58654 81922 58722 81978
rect 58778 81922 89318 81978
rect 89374 81922 89442 81978
rect 89498 81922 120038 81978
rect 120094 81922 120162 81978
rect 120218 81922 150758 81978
rect 150814 81922 150882 81978
rect 150938 81922 181478 81978
rect 181534 81922 181602 81978
rect 181658 81922 212198 81978
rect 212254 81922 212322 81978
rect 212378 81922 242918 81978
rect 242974 81922 243042 81978
rect 243098 81922 273638 81978
rect 273694 81922 273762 81978
rect 273818 81922 304358 81978
rect 304414 81922 304482 81978
rect 304538 81922 335078 81978
rect 335134 81922 335202 81978
rect 335258 81922 365798 81978
rect 365854 81922 365922 81978
rect 365978 81922 396518 81978
rect 396574 81922 396642 81978
rect 396698 81922 427238 81978
rect 427294 81922 427362 81978
rect 427418 81922 457958 81978
rect 458014 81922 458082 81978
rect 458138 81922 488678 81978
rect 488734 81922 488802 81978
rect 488858 81922 519398 81978
rect 519454 81922 519522 81978
rect 519578 81922 550118 81978
rect 550174 81922 550242 81978
rect 550298 81922 592914 81978
rect 592970 81922 593038 81978
rect 593094 81922 593162 81978
rect 593218 81922 593286 81978
rect 593342 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect -1916 81826 597980 81922
rect -1916 76350 597980 76446
rect -1916 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 5514 76350
rect 5570 76294 5638 76350
rect 5694 76294 5762 76350
rect 5818 76294 5886 76350
rect 5942 76294 12518 76350
rect 12574 76294 12642 76350
rect 12698 76294 43238 76350
rect 43294 76294 43362 76350
rect 43418 76294 73958 76350
rect 74014 76294 74082 76350
rect 74138 76294 104678 76350
rect 104734 76294 104802 76350
rect 104858 76294 135398 76350
rect 135454 76294 135522 76350
rect 135578 76294 166118 76350
rect 166174 76294 166242 76350
rect 166298 76294 196838 76350
rect 196894 76294 196962 76350
rect 197018 76294 227558 76350
rect 227614 76294 227682 76350
rect 227738 76294 258278 76350
rect 258334 76294 258402 76350
rect 258458 76294 288998 76350
rect 289054 76294 289122 76350
rect 289178 76294 319718 76350
rect 319774 76294 319842 76350
rect 319898 76294 350438 76350
rect 350494 76294 350562 76350
rect 350618 76294 381158 76350
rect 381214 76294 381282 76350
rect 381338 76294 411878 76350
rect 411934 76294 412002 76350
rect 412058 76294 442598 76350
rect 442654 76294 442722 76350
rect 442778 76294 473318 76350
rect 473374 76294 473442 76350
rect 473498 76294 504038 76350
rect 504094 76294 504162 76350
rect 504218 76294 534758 76350
rect 534814 76294 534882 76350
rect 534938 76294 565478 76350
rect 565534 76294 565602 76350
rect 565658 76294 589194 76350
rect 589250 76294 589318 76350
rect 589374 76294 589442 76350
rect 589498 76294 589566 76350
rect 589622 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597980 76350
rect -1916 76226 597980 76294
rect -1916 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 5514 76226
rect 5570 76170 5638 76226
rect 5694 76170 5762 76226
rect 5818 76170 5886 76226
rect 5942 76170 12518 76226
rect 12574 76170 12642 76226
rect 12698 76170 43238 76226
rect 43294 76170 43362 76226
rect 43418 76170 73958 76226
rect 74014 76170 74082 76226
rect 74138 76170 104678 76226
rect 104734 76170 104802 76226
rect 104858 76170 135398 76226
rect 135454 76170 135522 76226
rect 135578 76170 166118 76226
rect 166174 76170 166242 76226
rect 166298 76170 196838 76226
rect 196894 76170 196962 76226
rect 197018 76170 227558 76226
rect 227614 76170 227682 76226
rect 227738 76170 258278 76226
rect 258334 76170 258402 76226
rect 258458 76170 288998 76226
rect 289054 76170 289122 76226
rect 289178 76170 319718 76226
rect 319774 76170 319842 76226
rect 319898 76170 350438 76226
rect 350494 76170 350562 76226
rect 350618 76170 381158 76226
rect 381214 76170 381282 76226
rect 381338 76170 411878 76226
rect 411934 76170 412002 76226
rect 412058 76170 442598 76226
rect 442654 76170 442722 76226
rect 442778 76170 473318 76226
rect 473374 76170 473442 76226
rect 473498 76170 504038 76226
rect 504094 76170 504162 76226
rect 504218 76170 534758 76226
rect 534814 76170 534882 76226
rect 534938 76170 565478 76226
rect 565534 76170 565602 76226
rect 565658 76170 589194 76226
rect 589250 76170 589318 76226
rect 589374 76170 589442 76226
rect 589498 76170 589566 76226
rect 589622 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597980 76226
rect -1916 76102 597980 76170
rect -1916 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 5514 76102
rect 5570 76046 5638 76102
rect 5694 76046 5762 76102
rect 5818 76046 5886 76102
rect 5942 76046 12518 76102
rect 12574 76046 12642 76102
rect 12698 76046 43238 76102
rect 43294 76046 43362 76102
rect 43418 76046 73958 76102
rect 74014 76046 74082 76102
rect 74138 76046 104678 76102
rect 104734 76046 104802 76102
rect 104858 76046 135398 76102
rect 135454 76046 135522 76102
rect 135578 76046 166118 76102
rect 166174 76046 166242 76102
rect 166298 76046 196838 76102
rect 196894 76046 196962 76102
rect 197018 76046 227558 76102
rect 227614 76046 227682 76102
rect 227738 76046 258278 76102
rect 258334 76046 258402 76102
rect 258458 76046 288998 76102
rect 289054 76046 289122 76102
rect 289178 76046 319718 76102
rect 319774 76046 319842 76102
rect 319898 76046 350438 76102
rect 350494 76046 350562 76102
rect 350618 76046 381158 76102
rect 381214 76046 381282 76102
rect 381338 76046 411878 76102
rect 411934 76046 412002 76102
rect 412058 76046 442598 76102
rect 442654 76046 442722 76102
rect 442778 76046 473318 76102
rect 473374 76046 473442 76102
rect 473498 76046 504038 76102
rect 504094 76046 504162 76102
rect 504218 76046 534758 76102
rect 534814 76046 534882 76102
rect 534938 76046 565478 76102
rect 565534 76046 565602 76102
rect 565658 76046 589194 76102
rect 589250 76046 589318 76102
rect 589374 76046 589442 76102
rect 589498 76046 589566 76102
rect 589622 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597980 76102
rect -1916 75978 597980 76046
rect -1916 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 5514 75978
rect 5570 75922 5638 75978
rect 5694 75922 5762 75978
rect 5818 75922 5886 75978
rect 5942 75922 12518 75978
rect 12574 75922 12642 75978
rect 12698 75922 43238 75978
rect 43294 75922 43362 75978
rect 43418 75922 73958 75978
rect 74014 75922 74082 75978
rect 74138 75922 104678 75978
rect 104734 75922 104802 75978
rect 104858 75922 135398 75978
rect 135454 75922 135522 75978
rect 135578 75922 166118 75978
rect 166174 75922 166242 75978
rect 166298 75922 196838 75978
rect 196894 75922 196962 75978
rect 197018 75922 227558 75978
rect 227614 75922 227682 75978
rect 227738 75922 258278 75978
rect 258334 75922 258402 75978
rect 258458 75922 288998 75978
rect 289054 75922 289122 75978
rect 289178 75922 319718 75978
rect 319774 75922 319842 75978
rect 319898 75922 350438 75978
rect 350494 75922 350562 75978
rect 350618 75922 381158 75978
rect 381214 75922 381282 75978
rect 381338 75922 411878 75978
rect 411934 75922 412002 75978
rect 412058 75922 442598 75978
rect 442654 75922 442722 75978
rect 442778 75922 473318 75978
rect 473374 75922 473442 75978
rect 473498 75922 504038 75978
rect 504094 75922 504162 75978
rect 504218 75922 534758 75978
rect 534814 75922 534882 75978
rect 534938 75922 565478 75978
rect 565534 75922 565602 75978
rect 565658 75922 589194 75978
rect 589250 75922 589318 75978
rect 589374 75922 589442 75978
rect 589498 75922 589566 75978
rect 589622 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597980 75978
rect -1916 75826 597980 75922
rect -1916 64350 597980 64446
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 27878 64350
rect 27934 64294 28002 64350
rect 28058 64294 58598 64350
rect 58654 64294 58722 64350
rect 58778 64294 89318 64350
rect 89374 64294 89442 64350
rect 89498 64294 120038 64350
rect 120094 64294 120162 64350
rect 120218 64294 150758 64350
rect 150814 64294 150882 64350
rect 150938 64294 181478 64350
rect 181534 64294 181602 64350
rect 181658 64294 212198 64350
rect 212254 64294 212322 64350
rect 212378 64294 242918 64350
rect 242974 64294 243042 64350
rect 243098 64294 273638 64350
rect 273694 64294 273762 64350
rect 273818 64294 304358 64350
rect 304414 64294 304482 64350
rect 304538 64294 335078 64350
rect 335134 64294 335202 64350
rect 335258 64294 365798 64350
rect 365854 64294 365922 64350
rect 365978 64294 396518 64350
rect 396574 64294 396642 64350
rect 396698 64294 427238 64350
rect 427294 64294 427362 64350
rect 427418 64294 457958 64350
rect 458014 64294 458082 64350
rect 458138 64294 488678 64350
rect 488734 64294 488802 64350
rect 488858 64294 519398 64350
rect 519454 64294 519522 64350
rect 519578 64294 550118 64350
rect 550174 64294 550242 64350
rect 550298 64294 592914 64350
rect 592970 64294 593038 64350
rect 593094 64294 593162 64350
rect 593218 64294 593286 64350
rect 593342 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect -1916 64226 597980 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 27878 64226
rect 27934 64170 28002 64226
rect 28058 64170 58598 64226
rect 58654 64170 58722 64226
rect 58778 64170 89318 64226
rect 89374 64170 89442 64226
rect 89498 64170 120038 64226
rect 120094 64170 120162 64226
rect 120218 64170 150758 64226
rect 150814 64170 150882 64226
rect 150938 64170 181478 64226
rect 181534 64170 181602 64226
rect 181658 64170 212198 64226
rect 212254 64170 212322 64226
rect 212378 64170 242918 64226
rect 242974 64170 243042 64226
rect 243098 64170 273638 64226
rect 273694 64170 273762 64226
rect 273818 64170 304358 64226
rect 304414 64170 304482 64226
rect 304538 64170 335078 64226
rect 335134 64170 335202 64226
rect 335258 64170 365798 64226
rect 365854 64170 365922 64226
rect 365978 64170 396518 64226
rect 396574 64170 396642 64226
rect 396698 64170 427238 64226
rect 427294 64170 427362 64226
rect 427418 64170 457958 64226
rect 458014 64170 458082 64226
rect 458138 64170 488678 64226
rect 488734 64170 488802 64226
rect 488858 64170 519398 64226
rect 519454 64170 519522 64226
rect 519578 64170 550118 64226
rect 550174 64170 550242 64226
rect 550298 64170 592914 64226
rect 592970 64170 593038 64226
rect 593094 64170 593162 64226
rect 593218 64170 593286 64226
rect 593342 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect -1916 64102 597980 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 27878 64102
rect 27934 64046 28002 64102
rect 28058 64046 58598 64102
rect 58654 64046 58722 64102
rect 58778 64046 89318 64102
rect 89374 64046 89442 64102
rect 89498 64046 120038 64102
rect 120094 64046 120162 64102
rect 120218 64046 150758 64102
rect 150814 64046 150882 64102
rect 150938 64046 181478 64102
rect 181534 64046 181602 64102
rect 181658 64046 212198 64102
rect 212254 64046 212322 64102
rect 212378 64046 242918 64102
rect 242974 64046 243042 64102
rect 243098 64046 273638 64102
rect 273694 64046 273762 64102
rect 273818 64046 304358 64102
rect 304414 64046 304482 64102
rect 304538 64046 335078 64102
rect 335134 64046 335202 64102
rect 335258 64046 365798 64102
rect 365854 64046 365922 64102
rect 365978 64046 396518 64102
rect 396574 64046 396642 64102
rect 396698 64046 427238 64102
rect 427294 64046 427362 64102
rect 427418 64046 457958 64102
rect 458014 64046 458082 64102
rect 458138 64046 488678 64102
rect 488734 64046 488802 64102
rect 488858 64046 519398 64102
rect 519454 64046 519522 64102
rect 519578 64046 550118 64102
rect 550174 64046 550242 64102
rect 550298 64046 592914 64102
rect 592970 64046 593038 64102
rect 593094 64046 593162 64102
rect 593218 64046 593286 64102
rect 593342 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect -1916 63978 597980 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 27878 63978
rect 27934 63922 28002 63978
rect 28058 63922 58598 63978
rect 58654 63922 58722 63978
rect 58778 63922 89318 63978
rect 89374 63922 89442 63978
rect 89498 63922 120038 63978
rect 120094 63922 120162 63978
rect 120218 63922 150758 63978
rect 150814 63922 150882 63978
rect 150938 63922 181478 63978
rect 181534 63922 181602 63978
rect 181658 63922 212198 63978
rect 212254 63922 212322 63978
rect 212378 63922 242918 63978
rect 242974 63922 243042 63978
rect 243098 63922 273638 63978
rect 273694 63922 273762 63978
rect 273818 63922 304358 63978
rect 304414 63922 304482 63978
rect 304538 63922 335078 63978
rect 335134 63922 335202 63978
rect 335258 63922 365798 63978
rect 365854 63922 365922 63978
rect 365978 63922 396518 63978
rect 396574 63922 396642 63978
rect 396698 63922 427238 63978
rect 427294 63922 427362 63978
rect 427418 63922 457958 63978
rect 458014 63922 458082 63978
rect 458138 63922 488678 63978
rect 488734 63922 488802 63978
rect 488858 63922 519398 63978
rect 519454 63922 519522 63978
rect 519578 63922 550118 63978
rect 550174 63922 550242 63978
rect 550298 63922 592914 63978
rect 592970 63922 593038 63978
rect 593094 63922 593162 63978
rect 593218 63922 593286 63978
rect 593342 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect -1916 63826 597980 63922
rect -1916 58350 597980 58446
rect -1916 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 5514 58350
rect 5570 58294 5638 58350
rect 5694 58294 5762 58350
rect 5818 58294 5886 58350
rect 5942 58294 12518 58350
rect 12574 58294 12642 58350
rect 12698 58294 43238 58350
rect 43294 58294 43362 58350
rect 43418 58294 73958 58350
rect 74014 58294 74082 58350
rect 74138 58294 104678 58350
rect 104734 58294 104802 58350
rect 104858 58294 135398 58350
rect 135454 58294 135522 58350
rect 135578 58294 166118 58350
rect 166174 58294 166242 58350
rect 166298 58294 196838 58350
rect 196894 58294 196962 58350
rect 197018 58294 227558 58350
rect 227614 58294 227682 58350
rect 227738 58294 258278 58350
rect 258334 58294 258402 58350
rect 258458 58294 288998 58350
rect 289054 58294 289122 58350
rect 289178 58294 319718 58350
rect 319774 58294 319842 58350
rect 319898 58294 350438 58350
rect 350494 58294 350562 58350
rect 350618 58294 381158 58350
rect 381214 58294 381282 58350
rect 381338 58294 411878 58350
rect 411934 58294 412002 58350
rect 412058 58294 442598 58350
rect 442654 58294 442722 58350
rect 442778 58294 473318 58350
rect 473374 58294 473442 58350
rect 473498 58294 504038 58350
rect 504094 58294 504162 58350
rect 504218 58294 534758 58350
rect 534814 58294 534882 58350
rect 534938 58294 565478 58350
rect 565534 58294 565602 58350
rect 565658 58294 589194 58350
rect 589250 58294 589318 58350
rect 589374 58294 589442 58350
rect 589498 58294 589566 58350
rect 589622 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597980 58350
rect -1916 58226 597980 58294
rect -1916 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 5514 58226
rect 5570 58170 5638 58226
rect 5694 58170 5762 58226
rect 5818 58170 5886 58226
rect 5942 58170 12518 58226
rect 12574 58170 12642 58226
rect 12698 58170 43238 58226
rect 43294 58170 43362 58226
rect 43418 58170 73958 58226
rect 74014 58170 74082 58226
rect 74138 58170 104678 58226
rect 104734 58170 104802 58226
rect 104858 58170 135398 58226
rect 135454 58170 135522 58226
rect 135578 58170 166118 58226
rect 166174 58170 166242 58226
rect 166298 58170 196838 58226
rect 196894 58170 196962 58226
rect 197018 58170 227558 58226
rect 227614 58170 227682 58226
rect 227738 58170 258278 58226
rect 258334 58170 258402 58226
rect 258458 58170 288998 58226
rect 289054 58170 289122 58226
rect 289178 58170 319718 58226
rect 319774 58170 319842 58226
rect 319898 58170 350438 58226
rect 350494 58170 350562 58226
rect 350618 58170 381158 58226
rect 381214 58170 381282 58226
rect 381338 58170 411878 58226
rect 411934 58170 412002 58226
rect 412058 58170 442598 58226
rect 442654 58170 442722 58226
rect 442778 58170 473318 58226
rect 473374 58170 473442 58226
rect 473498 58170 504038 58226
rect 504094 58170 504162 58226
rect 504218 58170 534758 58226
rect 534814 58170 534882 58226
rect 534938 58170 565478 58226
rect 565534 58170 565602 58226
rect 565658 58170 589194 58226
rect 589250 58170 589318 58226
rect 589374 58170 589442 58226
rect 589498 58170 589566 58226
rect 589622 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597980 58226
rect -1916 58102 597980 58170
rect -1916 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 5514 58102
rect 5570 58046 5638 58102
rect 5694 58046 5762 58102
rect 5818 58046 5886 58102
rect 5942 58046 12518 58102
rect 12574 58046 12642 58102
rect 12698 58046 43238 58102
rect 43294 58046 43362 58102
rect 43418 58046 73958 58102
rect 74014 58046 74082 58102
rect 74138 58046 104678 58102
rect 104734 58046 104802 58102
rect 104858 58046 135398 58102
rect 135454 58046 135522 58102
rect 135578 58046 166118 58102
rect 166174 58046 166242 58102
rect 166298 58046 196838 58102
rect 196894 58046 196962 58102
rect 197018 58046 227558 58102
rect 227614 58046 227682 58102
rect 227738 58046 258278 58102
rect 258334 58046 258402 58102
rect 258458 58046 288998 58102
rect 289054 58046 289122 58102
rect 289178 58046 319718 58102
rect 319774 58046 319842 58102
rect 319898 58046 350438 58102
rect 350494 58046 350562 58102
rect 350618 58046 381158 58102
rect 381214 58046 381282 58102
rect 381338 58046 411878 58102
rect 411934 58046 412002 58102
rect 412058 58046 442598 58102
rect 442654 58046 442722 58102
rect 442778 58046 473318 58102
rect 473374 58046 473442 58102
rect 473498 58046 504038 58102
rect 504094 58046 504162 58102
rect 504218 58046 534758 58102
rect 534814 58046 534882 58102
rect 534938 58046 565478 58102
rect 565534 58046 565602 58102
rect 565658 58046 589194 58102
rect 589250 58046 589318 58102
rect 589374 58046 589442 58102
rect 589498 58046 589566 58102
rect 589622 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597980 58102
rect -1916 57978 597980 58046
rect -1916 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 5514 57978
rect 5570 57922 5638 57978
rect 5694 57922 5762 57978
rect 5818 57922 5886 57978
rect 5942 57922 12518 57978
rect 12574 57922 12642 57978
rect 12698 57922 43238 57978
rect 43294 57922 43362 57978
rect 43418 57922 73958 57978
rect 74014 57922 74082 57978
rect 74138 57922 104678 57978
rect 104734 57922 104802 57978
rect 104858 57922 135398 57978
rect 135454 57922 135522 57978
rect 135578 57922 166118 57978
rect 166174 57922 166242 57978
rect 166298 57922 196838 57978
rect 196894 57922 196962 57978
rect 197018 57922 227558 57978
rect 227614 57922 227682 57978
rect 227738 57922 258278 57978
rect 258334 57922 258402 57978
rect 258458 57922 288998 57978
rect 289054 57922 289122 57978
rect 289178 57922 319718 57978
rect 319774 57922 319842 57978
rect 319898 57922 350438 57978
rect 350494 57922 350562 57978
rect 350618 57922 381158 57978
rect 381214 57922 381282 57978
rect 381338 57922 411878 57978
rect 411934 57922 412002 57978
rect 412058 57922 442598 57978
rect 442654 57922 442722 57978
rect 442778 57922 473318 57978
rect 473374 57922 473442 57978
rect 473498 57922 504038 57978
rect 504094 57922 504162 57978
rect 504218 57922 534758 57978
rect 534814 57922 534882 57978
rect 534938 57922 565478 57978
rect 565534 57922 565602 57978
rect 565658 57922 589194 57978
rect 589250 57922 589318 57978
rect 589374 57922 589442 57978
rect 589498 57922 589566 57978
rect 589622 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597980 57978
rect -1916 57826 597980 57922
rect -1916 46350 597980 46446
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 27878 46350
rect 27934 46294 28002 46350
rect 28058 46294 58598 46350
rect 58654 46294 58722 46350
rect 58778 46294 89318 46350
rect 89374 46294 89442 46350
rect 89498 46294 120038 46350
rect 120094 46294 120162 46350
rect 120218 46294 150758 46350
rect 150814 46294 150882 46350
rect 150938 46294 181478 46350
rect 181534 46294 181602 46350
rect 181658 46294 212198 46350
rect 212254 46294 212322 46350
rect 212378 46294 242918 46350
rect 242974 46294 243042 46350
rect 243098 46294 273638 46350
rect 273694 46294 273762 46350
rect 273818 46294 304358 46350
rect 304414 46294 304482 46350
rect 304538 46294 335078 46350
rect 335134 46294 335202 46350
rect 335258 46294 365798 46350
rect 365854 46294 365922 46350
rect 365978 46294 396518 46350
rect 396574 46294 396642 46350
rect 396698 46294 427238 46350
rect 427294 46294 427362 46350
rect 427418 46294 457958 46350
rect 458014 46294 458082 46350
rect 458138 46294 488678 46350
rect 488734 46294 488802 46350
rect 488858 46294 519398 46350
rect 519454 46294 519522 46350
rect 519578 46294 550118 46350
rect 550174 46294 550242 46350
rect 550298 46294 592914 46350
rect 592970 46294 593038 46350
rect 593094 46294 593162 46350
rect 593218 46294 593286 46350
rect 593342 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect -1916 46226 597980 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 27878 46226
rect 27934 46170 28002 46226
rect 28058 46170 58598 46226
rect 58654 46170 58722 46226
rect 58778 46170 89318 46226
rect 89374 46170 89442 46226
rect 89498 46170 120038 46226
rect 120094 46170 120162 46226
rect 120218 46170 150758 46226
rect 150814 46170 150882 46226
rect 150938 46170 181478 46226
rect 181534 46170 181602 46226
rect 181658 46170 212198 46226
rect 212254 46170 212322 46226
rect 212378 46170 242918 46226
rect 242974 46170 243042 46226
rect 243098 46170 273638 46226
rect 273694 46170 273762 46226
rect 273818 46170 304358 46226
rect 304414 46170 304482 46226
rect 304538 46170 335078 46226
rect 335134 46170 335202 46226
rect 335258 46170 365798 46226
rect 365854 46170 365922 46226
rect 365978 46170 396518 46226
rect 396574 46170 396642 46226
rect 396698 46170 427238 46226
rect 427294 46170 427362 46226
rect 427418 46170 457958 46226
rect 458014 46170 458082 46226
rect 458138 46170 488678 46226
rect 488734 46170 488802 46226
rect 488858 46170 519398 46226
rect 519454 46170 519522 46226
rect 519578 46170 550118 46226
rect 550174 46170 550242 46226
rect 550298 46170 592914 46226
rect 592970 46170 593038 46226
rect 593094 46170 593162 46226
rect 593218 46170 593286 46226
rect 593342 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect -1916 46102 597980 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 27878 46102
rect 27934 46046 28002 46102
rect 28058 46046 58598 46102
rect 58654 46046 58722 46102
rect 58778 46046 89318 46102
rect 89374 46046 89442 46102
rect 89498 46046 120038 46102
rect 120094 46046 120162 46102
rect 120218 46046 150758 46102
rect 150814 46046 150882 46102
rect 150938 46046 181478 46102
rect 181534 46046 181602 46102
rect 181658 46046 212198 46102
rect 212254 46046 212322 46102
rect 212378 46046 242918 46102
rect 242974 46046 243042 46102
rect 243098 46046 273638 46102
rect 273694 46046 273762 46102
rect 273818 46046 304358 46102
rect 304414 46046 304482 46102
rect 304538 46046 335078 46102
rect 335134 46046 335202 46102
rect 335258 46046 365798 46102
rect 365854 46046 365922 46102
rect 365978 46046 396518 46102
rect 396574 46046 396642 46102
rect 396698 46046 427238 46102
rect 427294 46046 427362 46102
rect 427418 46046 457958 46102
rect 458014 46046 458082 46102
rect 458138 46046 488678 46102
rect 488734 46046 488802 46102
rect 488858 46046 519398 46102
rect 519454 46046 519522 46102
rect 519578 46046 550118 46102
rect 550174 46046 550242 46102
rect 550298 46046 592914 46102
rect 592970 46046 593038 46102
rect 593094 46046 593162 46102
rect 593218 46046 593286 46102
rect 593342 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect -1916 45978 597980 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 27878 45978
rect 27934 45922 28002 45978
rect 28058 45922 58598 45978
rect 58654 45922 58722 45978
rect 58778 45922 89318 45978
rect 89374 45922 89442 45978
rect 89498 45922 120038 45978
rect 120094 45922 120162 45978
rect 120218 45922 150758 45978
rect 150814 45922 150882 45978
rect 150938 45922 181478 45978
rect 181534 45922 181602 45978
rect 181658 45922 212198 45978
rect 212254 45922 212322 45978
rect 212378 45922 242918 45978
rect 242974 45922 243042 45978
rect 243098 45922 273638 45978
rect 273694 45922 273762 45978
rect 273818 45922 304358 45978
rect 304414 45922 304482 45978
rect 304538 45922 335078 45978
rect 335134 45922 335202 45978
rect 335258 45922 365798 45978
rect 365854 45922 365922 45978
rect 365978 45922 396518 45978
rect 396574 45922 396642 45978
rect 396698 45922 427238 45978
rect 427294 45922 427362 45978
rect 427418 45922 457958 45978
rect 458014 45922 458082 45978
rect 458138 45922 488678 45978
rect 488734 45922 488802 45978
rect 488858 45922 519398 45978
rect 519454 45922 519522 45978
rect 519578 45922 550118 45978
rect 550174 45922 550242 45978
rect 550298 45922 592914 45978
rect 592970 45922 593038 45978
rect 593094 45922 593162 45978
rect 593218 45922 593286 45978
rect 593342 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect -1916 45826 597980 45922
rect -1916 40350 597980 40446
rect -1916 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 5514 40350
rect 5570 40294 5638 40350
rect 5694 40294 5762 40350
rect 5818 40294 5886 40350
rect 5942 40294 12518 40350
rect 12574 40294 12642 40350
rect 12698 40294 43238 40350
rect 43294 40294 43362 40350
rect 43418 40294 73958 40350
rect 74014 40294 74082 40350
rect 74138 40294 104678 40350
rect 104734 40294 104802 40350
rect 104858 40294 135398 40350
rect 135454 40294 135522 40350
rect 135578 40294 166118 40350
rect 166174 40294 166242 40350
rect 166298 40294 196838 40350
rect 196894 40294 196962 40350
rect 197018 40294 227558 40350
rect 227614 40294 227682 40350
rect 227738 40294 258278 40350
rect 258334 40294 258402 40350
rect 258458 40294 288998 40350
rect 289054 40294 289122 40350
rect 289178 40294 319718 40350
rect 319774 40294 319842 40350
rect 319898 40294 350438 40350
rect 350494 40294 350562 40350
rect 350618 40294 381158 40350
rect 381214 40294 381282 40350
rect 381338 40294 411878 40350
rect 411934 40294 412002 40350
rect 412058 40294 442598 40350
rect 442654 40294 442722 40350
rect 442778 40294 473318 40350
rect 473374 40294 473442 40350
rect 473498 40294 504038 40350
rect 504094 40294 504162 40350
rect 504218 40294 534758 40350
rect 534814 40294 534882 40350
rect 534938 40294 565478 40350
rect 565534 40294 565602 40350
rect 565658 40294 589194 40350
rect 589250 40294 589318 40350
rect 589374 40294 589442 40350
rect 589498 40294 589566 40350
rect 589622 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597980 40350
rect -1916 40226 597980 40294
rect -1916 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 5514 40226
rect 5570 40170 5638 40226
rect 5694 40170 5762 40226
rect 5818 40170 5886 40226
rect 5942 40170 12518 40226
rect 12574 40170 12642 40226
rect 12698 40170 43238 40226
rect 43294 40170 43362 40226
rect 43418 40170 73958 40226
rect 74014 40170 74082 40226
rect 74138 40170 104678 40226
rect 104734 40170 104802 40226
rect 104858 40170 135398 40226
rect 135454 40170 135522 40226
rect 135578 40170 166118 40226
rect 166174 40170 166242 40226
rect 166298 40170 196838 40226
rect 196894 40170 196962 40226
rect 197018 40170 227558 40226
rect 227614 40170 227682 40226
rect 227738 40170 258278 40226
rect 258334 40170 258402 40226
rect 258458 40170 288998 40226
rect 289054 40170 289122 40226
rect 289178 40170 319718 40226
rect 319774 40170 319842 40226
rect 319898 40170 350438 40226
rect 350494 40170 350562 40226
rect 350618 40170 381158 40226
rect 381214 40170 381282 40226
rect 381338 40170 411878 40226
rect 411934 40170 412002 40226
rect 412058 40170 442598 40226
rect 442654 40170 442722 40226
rect 442778 40170 473318 40226
rect 473374 40170 473442 40226
rect 473498 40170 504038 40226
rect 504094 40170 504162 40226
rect 504218 40170 534758 40226
rect 534814 40170 534882 40226
rect 534938 40170 565478 40226
rect 565534 40170 565602 40226
rect 565658 40170 589194 40226
rect 589250 40170 589318 40226
rect 589374 40170 589442 40226
rect 589498 40170 589566 40226
rect 589622 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597980 40226
rect -1916 40102 597980 40170
rect -1916 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 5514 40102
rect 5570 40046 5638 40102
rect 5694 40046 5762 40102
rect 5818 40046 5886 40102
rect 5942 40046 12518 40102
rect 12574 40046 12642 40102
rect 12698 40046 43238 40102
rect 43294 40046 43362 40102
rect 43418 40046 73958 40102
rect 74014 40046 74082 40102
rect 74138 40046 104678 40102
rect 104734 40046 104802 40102
rect 104858 40046 135398 40102
rect 135454 40046 135522 40102
rect 135578 40046 166118 40102
rect 166174 40046 166242 40102
rect 166298 40046 196838 40102
rect 196894 40046 196962 40102
rect 197018 40046 227558 40102
rect 227614 40046 227682 40102
rect 227738 40046 258278 40102
rect 258334 40046 258402 40102
rect 258458 40046 288998 40102
rect 289054 40046 289122 40102
rect 289178 40046 319718 40102
rect 319774 40046 319842 40102
rect 319898 40046 350438 40102
rect 350494 40046 350562 40102
rect 350618 40046 381158 40102
rect 381214 40046 381282 40102
rect 381338 40046 411878 40102
rect 411934 40046 412002 40102
rect 412058 40046 442598 40102
rect 442654 40046 442722 40102
rect 442778 40046 473318 40102
rect 473374 40046 473442 40102
rect 473498 40046 504038 40102
rect 504094 40046 504162 40102
rect 504218 40046 534758 40102
rect 534814 40046 534882 40102
rect 534938 40046 565478 40102
rect 565534 40046 565602 40102
rect 565658 40046 589194 40102
rect 589250 40046 589318 40102
rect 589374 40046 589442 40102
rect 589498 40046 589566 40102
rect 589622 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597980 40102
rect -1916 39978 597980 40046
rect -1916 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 5514 39978
rect 5570 39922 5638 39978
rect 5694 39922 5762 39978
rect 5818 39922 5886 39978
rect 5942 39922 12518 39978
rect 12574 39922 12642 39978
rect 12698 39922 43238 39978
rect 43294 39922 43362 39978
rect 43418 39922 73958 39978
rect 74014 39922 74082 39978
rect 74138 39922 104678 39978
rect 104734 39922 104802 39978
rect 104858 39922 135398 39978
rect 135454 39922 135522 39978
rect 135578 39922 166118 39978
rect 166174 39922 166242 39978
rect 166298 39922 196838 39978
rect 196894 39922 196962 39978
rect 197018 39922 227558 39978
rect 227614 39922 227682 39978
rect 227738 39922 258278 39978
rect 258334 39922 258402 39978
rect 258458 39922 288998 39978
rect 289054 39922 289122 39978
rect 289178 39922 319718 39978
rect 319774 39922 319842 39978
rect 319898 39922 350438 39978
rect 350494 39922 350562 39978
rect 350618 39922 381158 39978
rect 381214 39922 381282 39978
rect 381338 39922 411878 39978
rect 411934 39922 412002 39978
rect 412058 39922 442598 39978
rect 442654 39922 442722 39978
rect 442778 39922 473318 39978
rect 473374 39922 473442 39978
rect 473498 39922 504038 39978
rect 504094 39922 504162 39978
rect 504218 39922 534758 39978
rect 534814 39922 534882 39978
rect 534938 39922 565478 39978
rect 565534 39922 565602 39978
rect 565658 39922 589194 39978
rect 589250 39922 589318 39978
rect 589374 39922 589442 39978
rect 589498 39922 589566 39978
rect 589622 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597980 39978
rect -1916 39826 597980 39922
rect -1916 28350 597980 28446
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 27878 28350
rect 27934 28294 28002 28350
rect 28058 28294 58598 28350
rect 58654 28294 58722 28350
rect 58778 28294 89318 28350
rect 89374 28294 89442 28350
rect 89498 28294 120038 28350
rect 120094 28294 120162 28350
rect 120218 28294 150758 28350
rect 150814 28294 150882 28350
rect 150938 28294 181478 28350
rect 181534 28294 181602 28350
rect 181658 28294 212198 28350
rect 212254 28294 212322 28350
rect 212378 28294 242918 28350
rect 242974 28294 243042 28350
rect 243098 28294 273638 28350
rect 273694 28294 273762 28350
rect 273818 28294 304358 28350
rect 304414 28294 304482 28350
rect 304538 28294 335078 28350
rect 335134 28294 335202 28350
rect 335258 28294 365798 28350
rect 365854 28294 365922 28350
rect 365978 28294 396518 28350
rect 396574 28294 396642 28350
rect 396698 28294 427238 28350
rect 427294 28294 427362 28350
rect 427418 28294 457958 28350
rect 458014 28294 458082 28350
rect 458138 28294 488678 28350
rect 488734 28294 488802 28350
rect 488858 28294 519398 28350
rect 519454 28294 519522 28350
rect 519578 28294 550118 28350
rect 550174 28294 550242 28350
rect 550298 28294 592914 28350
rect 592970 28294 593038 28350
rect 593094 28294 593162 28350
rect 593218 28294 593286 28350
rect 593342 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect -1916 28226 597980 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 27878 28226
rect 27934 28170 28002 28226
rect 28058 28170 58598 28226
rect 58654 28170 58722 28226
rect 58778 28170 89318 28226
rect 89374 28170 89442 28226
rect 89498 28170 120038 28226
rect 120094 28170 120162 28226
rect 120218 28170 150758 28226
rect 150814 28170 150882 28226
rect 150938 28170 181478 28226
rect 181534 28170 181602 28226
rect 181658 28170 212198 28226
rect 212254 28170 212322 28226
rect 212378 28170 242918 28226
rect 242974 28170 243042 28226
rect 243098 28170 273638 28226
rect 273694 28170 273762 28226
rect 273818 28170 304358 28226
rect 304414 28170 304482 28226
rect 304538 28170 335078 28226
rect 335134 28170 335202 28226
rect 335258 28170 365798 28226
rect 365854 28170 365922 28226
rect 365978 28170 396518 28226
rect 396574 28170 396642 28226
rect 396698 28170 427238 28226
rect 427294 28170 427362 28226
rect 427418 28170 457958 28226
rect 458014 28170 458082 28226
rect 458138 28170 488678 28226
rect 488734 28170 488802 28226
rect 488858 28170 519398 28226
rect 519454 28170 519522 28226
rect 519578 28170 550118 28226
rect 550174 28170 550242 28226
rect 550298 28170 592914 28226
rect 592970 28170 593038 28226
rect 593094 28170 593162 28226
rect 593218 28170 593286 28226
rect 593342 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect -1916 28102 597980 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 27878 28102
rect 27934 28046 28002 28102
rect 28058 28046 58598 28102
rect 58654 28046 58722 28102
rect 58778 28046 89318 28102
rect 89374 28046 89442 28102
rect 89498 28046 120038 28102
rect 120094 28046 120162 28102
rect 120218 28046 150758 28102
rect 150814 28046 150882 28102
rect 150938 28046 181478 28102
rect 181534 28046 181602 28102
rect 181658 28046 212198 28102
rect 212254 28046 212322 28102
rect 212378 28046 242918 28102
rect 242974 28046 243042 28102
rect 243098 28046 273638 28102
rect 273694 28046 273762 28102
rect 273818 28046 304358 28102
rect 304414 28046 304482 28102
rect 304538 28046 335078 28102
rect 335134 28046 335202 28102
rect 335258 28046 365798 28102
rect 365854 28046 365922 28102
rect 365978 28046 396518 28102
rect 396574 28046 396642 28102
rect 396698 28046 427238 28102
rect 427294 28046 427362 28102
rect 427418 28046 457958 28102
rect 458014 28046 458082 28102
rect 458138 28046 488678 28102
rect 488734 28046 488802 28102
rect 488858 28046 519398 28102
rect 519454 28046 519522 28102
rect 519578 28046 550118 28102
rect 550174 28046 550242 28102
rect 550298 28046 592914 28102
rect 592970 28046 593038 28102
rect 593094 28046 593162 28102
rect 593218 28046 593286 28102
rect 593342 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect -1916 27978 597980 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 27878 27978
rect 27934 27922 28002 27978
rect 28058 27922 58598 27978
rect 58654 27922 58722 27978
rect 58778 27922 89318 27978
rect 89374 27922 89442 27978
rect 89498 27922 120038 27978
rect 120094 27922 120162 27978
rect 120218 27922 150758 27978
rect 150814 27922 150882 27978
rect 150938 27922 181478 27978
rect 181534 27922 181602 27978
rect 181658 27922 212198 27978
rect 212254 27922 212322 27978
rect 212378 27922 242918 27978
rect 242974 27922 243042 27978
rect 243098 27922 273638 27978
rect 273694 27922 273762 27978
rect 273818 27922 304358 27978
rect 304414 27922 304482 27978
rect 304538 27922 335078 27978
rect 335134 27922 335202 27978
rect 335258 27922 365798 27978
rect 365854 27922 365922 27978
rect 365978 27922 396518 27978
rect 396574 27922 396642 27978
rect 396698 27922 427238 27978
rect 427294 27922 427362 27978
rect 427418 27922 457958 27978
rect 458014 27922 458082 27978
rect 458138 27922 488678 27978
rect 488734 27922 488802 27978
rect 488858 27922 519398 27978
rect 519454 27922 519522 27978
rect 519578 27922 550118 27978
rect 550174 27922 550242 27978
rect 550298 27922 592914 27978
rect 592970 27922 593038 27978
rect 593094 27922 593162 27978
rect 593218 27922 593286 27978
rect 593342 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect -1916 27826 597980 27922
rect -1916 22350 597980 22446
rect -1916 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 5514 22350
rect 5570 22294 5638 22350
rect 5694 22294 5762 22350
rect 5818 22294 5886 22350
rect 5942 22294 12518 22350
rect 12574 22294 12642 22350
rect 12698 22294 43238 22350
rect 43294 22294 43362 22350
rect 43418 22294 73958 22350
rect 74014 22294 74082 22350
rect 74138 22294 104678 22350
rect 104734 22294 104802 22350
rect 104858 22294 135398 22350
rect 135454 22294 135522 22350
rect 135578 22294 166118 22350
rect 166174 22294 166242 22350
rect 166298 22294 196838 22350
rect 196894 22294 196962 22350
rect 197018 22294 227558 22350
rect 227614 22294 227682 22350
rect 227738 22294 258278 22350
rect 258334 22294 258402 22350
rect 258458 22294 288998 22350
rect 289054 22294 289122 22350
rect 289178 22294 319718 22350
rect 319774 22294 319842 22350
rect 319898 22294 350438 22350
rect 350494 22294 350562 22350
rect 350618 22294 381158 22350
rect 381214 22294 381282 22350
rect 381338 22294 411878 22350
rect 411934 22294 412002 22350
rect 412058 22294 442598 22350
rect 442654 22294 442722 22350
rect 442778 22294 473318 22350
rect 473374 22294 473442 22350
rect 473498 22294 504038 22350
rect 504094 22294 504162 22350
rect 504218 22294 534758 22350
rect 534814 22294 534882 22350
rect 534938 22294 565478 22350
rect 565534 22294 565602 22350
rect 565658 22294 589194 22350
rect 589250 22294 589318 22350
rect 589374 22294 589442 22350
rect 589498 22294 589566 22350
rect 589622 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597980 22350
rect -1916 22226 597980 22294
rect -1916 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 5514 22226
rect 5570 22170 5638 22226
rect 5694 22170 5762 22226
rect 5818 22170 5886 22226
rect 5942 22170 12518 22226
rect 12574 22170 12642 22226
rect 12698 22170 43238 22226
rect 43294 22170 43362 22226
rect 43418 22170 73958 22226
rect 74014 22170 74082 22226
rect 74138 22170 104678 22226
rect 104734 22170 104802 22226
rect 104858 22170 135398 22226
rect 135454 22170 135522 22226
rect 135578 22170 166118 22226
rect 166174 22170 166242 22226
rect 166298 22170 196838 22226
rect 196894 22170 196962 22226
rect 197018 22170 227558 22226
rect 227614 22170 227682 22226
rect 227738 22170 258278 22226
rect 258334 22170 258402 22226
rect 258458 22170 288998 22226
rect 289054 22170 289122 22226
rect 289178 22170 319718 22226
rect 319774 22170 319842 22226
rect 319898 22170 350438 22226
rect 350494 22170 350562 22226
rect 350618 22170 381158 22226
rect 381214 22170 381282 22226
rect 381338 22170 411878 22226
rect 411934 22170 412002 22226
rect 412058 22170 442598 22226
rect 442654 22170 442722 22226
rect 442778 22170 473318 22226
rect 473374 22170 473442 22226
rect 473498 22170 504038 22226
rect 504094 22170 504162 22226
rect 504218 22170 534758 22226
rect 534814 22170 534882 22226
rect 534938 22170 565478 22226
rect 565534 22170 565602 22226
rect 565658 22170 589194 22226
rect 589250 22170 589318 22226
rect 589374 22170 589442 22226
rect 589498 22170 589566 22226
rect 589622 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597980 22226
rect -1916 22102 597980 22170
rect -1916 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 5514 22102
rect 5570 22046 5638 22102
rect 5694 22046 5762 22102
rect 5818 22046 5886 22102
rect 5942 22046 12518 22102
rect 12574 22046 12642 22102
rect 12698 22046 43238 22102
rect 43294 22046 43362 22102
rect 43418 22046 73958 22102
rect 74014 22046 74082 22102
rect 74138 22046 104678 22102
rect 104734 22046 104802 22102
rect 104858 22046 135398 22102
rect 135454 22046 135522 22102
rect 135578 22046 166118 22102
rect 166174 22046 166242 22102
rect 166298 22046 196838 22102
rect 196894 22046 196962 22102
rect 197018 22046 227558 22102
rect 227614 22046 227682 22102
rect 227738 22046 258278 22102
rect 258334 22046 258402 22102
rect 258458 22046 288998 22102
rect 289054 22046 289122 22102
rect 289178 22046 319718 22102
rect 319774 22046 319842 22102
rect 319898 22046 350438 22102
rect 350494 22046 350562 22102
rect 350618 22046 381158 22102
rect 381214 22046 381282 22102
rect 381338 22046 411878 22102
rect 411934 22046 412002 22102
rect 412058 22046 442598 22102
rect 442654 22046 442722 22102
rect 442778 22046 473318 22102
rect 473374 22046 473442 22102
rect 473498 22046 504038 22102
rect 504094 22046 504162 22102
rect 504218 22046 534758 22102
rect 534814 22046 534882 22102
rect 534938 22046 565478 22102
rect 565534 22046 565602 22102
rect 565658 22046 589194 22102
rect 589250 22046 589318 22102
rect 589374 22046 589442 22102
rect 589498 22046 589566 22102
rect 589622 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597980 22102
rect -1916 21978 597980 22046
rect -1916 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 5514 21978
rect 5570 21922 5638 21978
rect 5694 21922 5762 21978
rect 5818 21922 5886 21978
rect 5942 21922 12518 21978
rect 12574 21922 12642 21978
rect 12698 21922 43238 21978
rect 43294 21922 43362 21978
rect 43418 21922 73958 21978
rect 74014 21922 74082 21978
rect 74138 21922 104678 21978
rect 104734 21922 104802 21978
rect 104858 21922 135398 21978
rect 135454 21922 135522 21978
rect 135578 21922 166118 21978
rect 166174 21922 166242 21978
rect 166298 21922 196838 21978
rect 196894 21922 196962 21978
rect 197018 21922 227558 21978
rect 227614 21922 227682 21978
rect 227738 21922 258278 21978
rect 258334 21922 258402 21978
rect 258458 21922 288998 21978
rect 289054 21922 289122 21978
rect 289178 21922 319718 21978
rect 319774 21922 319842 21978
rect 319898 21922 350438 21978
rect 350494 21922 350562 21978
rect 350618 21922 381158 21978
rect 381214 21922 381282 21978
rect 381338 21922 411878 21978
rect 411934 21922 412002 21978
rect 412058 21922 442598 21978
rect 442654 21922 442722 21978
rect 442778 21922 473318 21978
rect 473374 21922 473442 21978
rect 473498 21922 504038 21978
rect 504094 21922 504162 21978
rect 504218 21922 534758 21978
rect 534814 21922 534882 21978
rect 534938 21922 565478 21978
rect 565534 21922 565602 21978
rect 565658 21922 589194 21978
rect 589250 21922 589318 21978
rect 589374 21922 589442 21978
rect 589498 21922 589566 21978
rect 589622 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597980 21978
rect -1916 21826 597980 21922
rect -1916 10350 597980 10446
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 592914 10350
rect 592970 10294 593038 10350
rect 593094 10294 593162 10350
rect 593218 10294 593286 10350
rect 593342 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect -1916 10226 597980 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 592914 10226
rect 592970 10170 593038 10226
rect 593094 10170 593162 10226
rect 593218 10170 593286 10226
rect 593342 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect -1916 10102 597980 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 592914 10102
rect 592970 10046 593038 10102
rect 593094 10046 593162 10102
rect 593218 10046 593286 10102
rect 593342 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect -1916 9978 597980 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 592914 9978
rect 592970 9922 593038 9978
rect 593094 9922 593162 9978
rect 593218 9922 593286 9978
rect 593342 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect -1916 9826 597980 9922
rect 557436 4978 576900 4994
rect 557436 4922 557452 4978
rect 557508 4922 576828 4978
rect 576884 4922 576900 4978
rect 557436 4906 576900 4922
rect 561020 4798 580708 4814
rect 561020 4742 561036 4798
rect 561092 4742 580636 4798
rect 580692 4742 580708 4798
rect 561020 4726 580708 4742
rect -1916 4350 597980 4446
rect -1916 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 5514 4350
rect 5570 4294 5638 4350
rect 5694 4294 5762 4350
rect 5818 4294 5886 4350
rect 5942 4294 36234 4350
rect 36290 4294 36358 4350
rect 36414 4294 36482 4350
rect 36538 4294 36606 4350
rect 36662 4294 66954 4350
rect 67010 4294 67078 4350
rect 67134 4294 67202 4350
rect 67258 4294 67326 4350
rect 67382 4294 97674 4350
rect 97730 4294 97798 4350
rect 97854 4294 97922 4350
rect 97978 4294 98046 4350
rect 98102 4294 128394 4350
rect 128450 4294 128518 4350
rect 128574 4294 128642 4350
rect 128698 4294 128766 4350
rect 128822 4294 159114 4350
rect 159170 4294 159238 4350
rect 159294 4294 159362 4350
rect 159418 4294 159486 4350
rect 159542 4294 189834 4350
rect 189890 4294 189958 4350
rect 190014 4294 190082 4350
rect 190138 4294 190206 4350
rect 190262 4294 220554 4350
rect 220610 4294 220678 4350
rect 220734 4294 220802 4350
rect 220858 4294 220926 4350
rect 220982 4294 251274 4350
rect 251330 4294 251398 4350
rect 251454 4294 251522 4350
rect 251578 4294 251646 4350
rect 251702 4294 281994 4350
rect 282050 4294 282118 4350
rect 282174 4294 282242 4350
rect 282298 4294 282366 4350
rect 282422 4294 312714 4350
rect 312770 4294 312838 4350
rect 312894 4294 312962 4350
rect 313018 4294 313086 4350
rect 313142 4294 343434 4350
rect 343490 4294 343558 4350
rect 343614 4294 343682 4350
rect 343738 4294 343806 4350
rect 343862 4294 374154 4350
rect 374210 4294 374278 4350
rect 374334 4294 374402 4350
rect 374458 4294 374526 4350
rect 374582 4294 404874 4350
rect 404930 4294 404998 4350
rect 405054 4294 405122 4350
rect 405178 4294 405246 4350
rect 405302 4294 435594 4350
rect 435650 4294 435718 4350
rect 435774 4294 435842 4350
rect 435898 4294 435966 4350
rect 436022 4294 466314 4350
rect 466370 4294 466438 4350
rect 466494 4294 466562 4350
rect 466618 4294 466686 4350
rect 466742 4294 497034 4350
rect 497090 4294 497158 4350
rect 497214 4294 497282 4350
rect 497338 4294 497406 4350
rect 497462 4294 527754 4350
rect 527810 4294 527878 4350
rect 527934 4294 528002 4350
rect 528058 4294 528126 4350
rect 528182 4294 558474 4350
rect 558530 4294 558598 4350
rect 558654 4294 558722 4350
rect 558778 4294 558846 4350
rect 558902 4294 589194 4350
rect 589250 4294 589318 4350
rect 589374 4294 589442 4350
rect 589498 4294 589566 4350
rect 589622 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597980 4350
rect -1916 4226 597980 4294
rect -1916 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 5514 4226
rect 5570 4170 5638 4226
rect 5694 4170 5762 4226
rect 5818 4170 5886 4226
rect 5942 4170 36234 4226
rect 36290 4170 36358 4226
rect 36414 4170 36482 4226
rect 36538 4170 36606 4226
rect 36662 4170 66954 4226
rect 67010 4170 67078 4226
rect 67134 4170 67202 4226
rect 67258 4170 67326 4226
rect 67382 4170 97674 4226
rect 97730 4170 97798 4226
rect 97854 4170 97922 4226
rect 97978 4170 98046 4226
rect 98102 4170 128394 4226
rect 128450 4170 128518 4226
rect 128574 4170 128642 4226
rect 128698 4170 128766 4226
rect 128822 4170 159114 4226
rect 159170 4170 159238 4226
rect 159294 4170 159362 4226
rect 159418 4170 159486 4226
rect 159542 4170 189834 4226
rect 189890 4170 189958 4226
rect 190014 4170 190082 4226
rect 190138 4170 190206 4226
rect 190262 4170 220554 4226
rect 220610 4170 220678 4226
rect 220734 4170 220802 4226
rect 220858 4170 220926 4226
rect 220982 4170 251274 4226
rect 251330 4170 251398 4226
rect 251454 4170 251522 4226
rect 251578 4170 251646 4226
rect 251702 4170 281994 4226
rect 282050 4170 282118 4226
rect 282174 4170 282242 4226
rect 282298 4170 282366 4226
rect 282422 4170 312714 4226
rect 312770 4170 312838 4226
rect 312894 4170 312962 4226
rect 313018 4170 313086 4226
rect 313142 4170 343434 4226
rect 343490 4170 343558 4226
rect 343614 4170 343682 4226
rect 343738 4170 343806 4226
rect 343862 4170 374154 4226
rect 374210 4170 374278 4226
rect 374334 4170 374402 4226
rect 374458 4170 374526 4226
rect 374582 4170 404874 4226
rect 404930 4170 404998 4226
rect 405054 4170 405122 4226
rect 405178 4170 405246 4226
rect 405302 4170 435594 4226
rect 435650 4170 435718 4226
rect 435774 4170 435842 4226
rect 435898 4170 435966 4226
rect 436022 4170 466314 4226
rect 466370 4170 466438 4226
rect 466494 4170 466562 4226
rect 466618 4170 466686 4226
rect 466742 4170 497034 4226
rect 497090 4170 497158 4226
rect 497214 4170 497282 4226
rect 497338 4170 497406 4226
rect 497462 4170 527754 4226
rect 527810 4170 527878 4226
rect 527934 4170 528002 4226
rect 528058 4170 528126 4226
rect 528182 4170 558474 4226
rect 558530 4170 558598 4226
rect 558654 4170 558722 4226
rect 558778 4170 558846 4226
rect 558902 4170 589194 4226
rect 589250 4170 589318 4226
rect 589374 4170 589442 4226
rect 589498 4170 589566 4226
rect 589622 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597980 4226
rect -1916 4102 597980 4170
rect -1916 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 5514 4102
rect 5570 4046 5638 4102
rect 5694 4046 5762 4102
rect 5818 4046 5886 4102
rect 5942 4046 36234 4102
rect 36290 4046 36358 4102
rect 36414 4046 36482 4102
rect 36538 4046 36606 4102
rect 36662 4046 66954 4102
rect 67010 4046 67078 4102
rect 67134 4046 67202 4102
rect 67258 4046 67326 4102
rect 67382 4046 97674 4102
rect 97730 4046 97798 4102
rect 97854 4046 97922 4102
rect 97978 4046 98046 4102
rect 98102 4046 128394 4102
rect 128450 4046 128518 4102
rect 128574 4046 128642 4102
rect 128698 4046 128766 4102
rect 128822 4046 159114 4102
rect 159170 4046 159238 4102
rect 159294 4046 159362 4102
rect 159418 4046 159486 4102
rect 159542 4046 189834 4102
rect 189890 4046 189958 4102
rect 190014 4046 190082 4102
rect 190138 4046 190206 4102
rect 190262 4046 220554 4102
rect 220610 4046 220678 4102
rect 220734 4046 220802 4102
rect 220858 4046 220926 4102
rect 220982 4046 251274 4102
rect 251330 4046 251398 4102
rect 251454 4046 251522 4102
rect 251578 4046 251646 4102
rect 251702 4046 281994 4102
rect 282050 4046 282118 4102
rect 282174 4046 282242 4102
rect 282298 4046 282366 4102
rect 282422 4046 312714 4102
rect 312770 4046 312838 4102
rect 312894 4046 312962 4102
rect 313018 4046 313086 4102
rect 313142 4046 343434 4102
rect 343490 4046 343558 4102
rect 343614 4046 343682 4102
rect 343738 4046 343806 4102
rect 343862 4046 374154 4102
rect 374210 4046 374278 4102
rect 374334 4046 374402 4102
rect 374458 4046 374526 4102
rect 374582 4046 404874 4102
rect 404930 4046 404998 4102
rect 405054 4046 405122 4102
rect 405178 4046 405246 4102
rect 405302 4046 435594 4102
rect 435650 4046 435718 4102
rect 435774 4046 435842 4102
rect 435898 4046 435966 4102
rect 436022 4046 466314 4102
rect 466370 4046 466438 4102
rect 466494 4046 466562 4102
rect 466618 4046 466686 4102
rect 466742 4046 497034 4102
rect 497090 4046 497158 4102
rect 497214 4046 497282 4102
rect 497338 4046 497406 4102
rect 497462 4046 527754 4102
rect 527810 4046 527878 4102
rect 527934 4046 528002 4102
rect 528058 4046 528126 4102
rect 528182 4046 558474 4102
rect 558530 4046 558598 4102
rect 558654 4046 558722 4102
rect 558778 4046 558846 4102
rect 558902 4046 589194 4102
rect 589250 4046 589318 4102
rect 589374 4046 589442 4102
rect 589498 4046 589566 4102
rect 589622 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597980 4102
rect -1916 3978 597980 4046
rect -1916 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 5514 3978
rect 5570 3922 5638 3978
rect 5694 3922 5762 3978
rect 5818 3922 5886 3978
rect 5942 3922 36234 3978
rect 36290 3922 36358 3978
rect 36414 3922 36482 3978
rect 36538 3922 36606 3978
rect 36662 3922 66954 3978
rect 67010 3922 67078 3978
rect 67134 3922 67202 3978
rect 67258 3922 67326 3978
rect 67382 3922 97674 3978
rect 97730 3922 97798 3978
rect 97854 3922 97922 3978
rect 97978 3922 98046 3978
rect 98102 3922 128394 3978
rect 128450 3922 128518 3978
rect 128574 3922 128642 3978
rect 128698 3922 128766 3978
rect 128822 3922 159114 3978
rect 159170 3922 159238 3978
rect 159294 3922 159362 3978
rect 159418 3922 159486 3978
rect 159542 3922 189834 3978
rect 189890 3922 189958 3978
rect 190014 3922 190082 3978
rect 190138 3922 190206 3978
rect 190262 3922 220554 3978
rect 220610 3922 220678 3978
rect 220734 3922 220802 3978
rect 220858 3922 220926 3978
rect 220982 3922 251274 3978
rect 251330 3922 251398 3978
rect 251454 3922 251522 3978
rect 251578 3922 251646 3978
rect 251702 3922 281994 3978
rect 282050 3922 282118 3978
rect 282174 3922 282242 3978
rect 282298 3922 282366 3978
rect 282422 3922 312714 3978
rect 312770 3922 312838 3978
rect 312894 3922 312962 3978
rect 313018 3922 313086 3978
rect 313142 3922 343434 3978
rect 343490 3922 343558 3978
rect 343614 3922 343682 3978
rect 343738 3922 343806 3978
rect 343862 3922 374154 3978
rect 374210 3922 374278 3978
rect 374334 3922 374402 3978
rect 374458 3922 374526 3978
rect 374582 3922 404874 3978
rect 404930 3922 404998 3978
rect 405054 3922 405122 3978
rect 405178 3922 405246 3978
rect 405302 3922 435594 3978
rect 435650 3922 435718 3978
rect 435774 3922 435842 3978
rect 435898 3922 435966 3978
rect 436022 3922 466314 3978
rect 466370 3922 466438 3978
rect 466494 3922 466562 3978
rect 466618 3922 466686 3978
rect 466742 3922 497034 3978
rect 497090 3922 497158 3978
rect 497214 3922 497282 3978
rect 497338 3922 497406 3978
rect 497462 3922 527754 3978
rect 527810 3922 527878 3978
rect 527934 3922 528002 3978
rect 528058 3922 528126 3978
rect 528182 3922 558474 3978
rect 558530 3922 558598 3978
rect 558654 3922 558722 3978
rect 558778 3922 558846 3978
rect 558902 3922 589194 3978
rect 589250 3922 589318 3978
rect 589374 3922 589442 3978
rect 589498 3922 589566 3978
rect 589622 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597980 3978
rect -1916 3826 597980 3922
rect -956 -160 597020 -64
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 5514 -160
rect 5570 -216 5638 -160
rect 5694 -216 5762 -160
rect 5818 -216 5886 -160
rect 5942 -216 36234 -160
rect 36290 -216 36358 -160
rect 36414 -216 36482 -160
rect 36538 -216 36606 -160
rect 36662 -216 66954 -160
rect 67010 -216 67078 -160
rect 67134 -216 67202 -160
rect 67258 -216 67326 -160
rect 67382 -216 97674 -160
rect 97730 -216 97798 -160
rect 97854 -216 97922 -160
rect 97978 -216 98046 -160
rect 98102 -216 128394 -160
rect 128450 -216 128518 -160
rect 128574 -216 128642 -160
rect 128698 -216 128766 -160
rect 128822 -216 159114 -160
rect 159170 -216 159238 -160
rect 159294 -216 159362 -160
rect 159418 -216 159486 -160
rect 159542 -216 189834 -160
rect 189890 -216 189958 -160
rect 190014 -216 190082 -160
rect 190138 -216 190206 -160
rect 190262 -216 220554 -160
rect 220610 -216 220678 -160
rect 220734 -216 220802 -160
rect 220858 -216 220926 -160
rect 220982 -216 251274 -160
rect 251330 -216 251398 -160
rect 251454 -216 251522 -160
rect 251578 -216 251646 -160
rect 251702 -216 281994 -160
rect 282050 -216 282118 -160
rect 282174 -216 282242 -160
rect 282298 -216 282366 -160
rect 282422 -216 312714 -160
rect 312770 -216 312838 -160
rect 312894 -216 312962 -160
rect 313018 -216 313086 -160
rect 313142 -216 343434 -160
rect 343490 -216 343558 -160
rect 343614 -216 343682 -160
rect 343738 -216 343806 -160
rect 343862 -216 374154 -160
rect 374210 -216 374278 -160
rect 374334 -216 374402 -160
rect 374458 -216 374526 -160
rect 374582 -216 404874 -160
rect 404930 -216 404998 -160
rect 405054 -216 405122 -160
rect 405178 -216 405246 -160
rect 405302 -216 435594 -160
rect 435650 -216 435718 -160
rect 435774 -216 435842 -160
rect 435898 -216 435966 -160
rect 436022 -216 466314 -160
rect 466370 -216 466438 -160
rect 466494 -216 466562 -160
rect 466618 -216 466686 -160
rect 466742 -216 497034 -160
rect 497090 -216 497158 -160
rect 497214 -216 497282 -160
rect 497338 -216 497406 -160
rect 497462 -216 527754 -160
rect 527810 -216 527878 -160
rect 527934 -216 528002 -160
rect 528058 -216 528126 -160
rect 528182 -216 558474 -160
rect 558530 -216 558598 -160
rect 558654 -216 558722 -160
rect 558778 -216 558846 -160
rect 558902 -216 589194 -160
rect 589250 -216 589318 -160
rect 589374 -216 589442 -160
rect 589498 -216 589566 -160
rect 589622 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect -956 -284 597020 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 5514 -284
rect 5570 -340 5638 -284
rect 5694 -340 5762 -284
rect 5818 -340 5886 -284
rect 5942 -340 36234 -284
rect 36290 -340 36358 -284
rect 36414 -340 36482 -284
rect 36538 -340 36606 -284
rect 36662 -340 66954 -284
rect 67010 -340 67078 -284
rect 67134 -340 67202 -284
rect 67258 -340 67326 -284
rect 67382 -340 97674 -284
rect 97730 -340 97798 -284
rect 97854 -340 97922 -284
rect 97978 -340 98046 -284
rect 98102 -340 128394 -284
rect 128450 -340 128518 -284
rect 128574 -340 128642 -284
rect 128698 -340 128766 -284
rect 128822 -340 159114 -284
rect 159170 -340 159238 -284
rect 159294 -340 159362 -284
rect 159418 -340 159486 -284
rect 159542 -340 189834 -284
rect 189890 -340 189958 -284
rect 190014 -340 190082 -284
rect 190138 -340 190206 -284
rect 190262 -340 220554 -284
rect 220610 -340 220678 -284
rect 220734 -340 220802 -284
rect 220858 -340 220926 -284
rect 220982 -340 251274 -284
rect 251330 -340 251398 -284
rect 251454 -340 251522 -284
rect 251578 -340 251646 -284
rect 251702 -340 281994 -284
rect 282050 -340 282118 -284
rect 282174 -340 282242 -284
rect 282298 -340 282366 -284
rect 282422 -340 312714 -284
rect 312770 -340 312838 -284
rect 312894 -340 312962 -284
rect 313018 -340 313086 -284
rect 313142 -340 343434 -284
rect 343490 -340 343558 -284
rect 343614 -340 343682 -284
rect 343738 -340 343806 -284
rect 343862 -340 374154 -284
rect 374210 -340 374278 -284
rect 374334 -340 374402 -284
rect 374458 -340 374526 -284
rect 374582 -340 404874 -284
rect 404930 -340 404998 -284
rect 405054 -340 405122 -284
rect 405178 -340 405246 -284
rect 405302 -340 435594 -284
rect 435650 -340 435718 -284
rect 435774 -340 435842 -284
rect 435898 -340 435966 -284
rect 436022 -340 466314 -284
rect 466370 -340 466438 -284
rect 466494 -340 466562 -284
rect 466618 -340 466686 -284
rect 466742 -340 497034 -284
rect 497090 -340 497158 -284
rect 497214 -340 497282 -284
rect 497338 -340 497406 -284
rect 497462 -340 527754 -284
rect 527810 -340 527878 -284
rect 527934 -340 528002 -284
rect 528058 -340 528126 -284
rect 528182 -340 558474 -284
rect 558530 -340 558598 -284
rect 558654 -340 558722 -284
rect 558778 -340 558846 -284
rect 558902 -340 589194 -284
rect 589250 -340 589318 -284
rect 589374 -340 589442 -284
rect 589498 -340 589566 -284
rect 589622 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect -956 -408 597020 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 5514 -408
rect 5570 -464 5638 -408
rect 5694 -464 5762 -408
rect 5818 -464 5886 -408
rect 5942 -464 36234 -408
rect 36290 -464 36358 -408
rect 36414 -464 36482 -408
rect 36538 -464 36606 -408
rect 36662 -464 66954 -408
rect 67010 -464 67078 -408
rect 67134 -464 67202 -408
rect 67258 -464 67326 -408
rect 67382 -464 97674 -408
rect 97730 -464 97798 -408
rect 97854 -464 97922 -408
rect 97978 -464 98046 -408
rect 98102 -464 128394 -408
rect 128450 -464 128518 -408
rect 128574 -464 128642 -408
rect 128698 -464 128766 -408
rect 128822 -464 159114 -408
rect 159170 -464 159238 -408
rect 159294 -464 159362 -408
rect 159418 -464 159486 -408
rect 159542 -464 189834 -408
rect 189890 -464 189958 -408
rect 190014 -464 190082 -408
rect 190138 -464 190206 -408
rect 190262 -464 220554 -408
rect 220610 -464 220678 -408
rect 220734 -464 220802 -408
rect 220858 -464 220926 -408
rect 220982 -464 251274 -408
rect 251330 -464 251398 -408
rect 251454 -464 251522 -408
rect 251578 -464 251646 -408
rect 251702 -464 281994 -408
rect 282050 -464 282118 -408
rect 282174 -464 282242 -408
rect 282298 -464 282366 -408
rect 282422 -464 312714 -408
rect 312770 -464 312838 -408
rect 312894 -464 312962 -408
rect 313018 -464 313086 -408
rect 313142 -464 343434 -408
rect 343490 -464 343558 -408
rect 343614 -464 343682 -408
rect 343738 -464 343806 -408
rect 343862 -464 374154 -408
rect 374210 -464 374278 -408
rect 374334 -464 374402 -408
rect 374458 -464 374526 -408
rect 374582 -464 404874 -408
rect 404930 -464 404998 -408
rect 405054 -464 405122 -408
rect 405178 -464 405246 -408
rect 405302 -464 435594 -408
rect 435650 -464 435718 -408
rect 435774 -464 435842 -408
rect 435898 -464 435966 -408
rect 436022 -464 466314 -408
rect 466370 -464 466438 -408
rect 466494 -464 466562 -408
rect 466618 -464 466686 -408
rect 466742 -464 497034 -408
rect 497090 -464 497158 -408
rect 497214 -464 497282 -408
rect 497338 -464 497406 -408
rect 497462 -464 527754 -408
rect 527810 -464 527878 -408
rect 527934 -464 528002 -408
rect 528058 -464 528126 -408
rect 528182 -464 558474 -408
rect 558530 -464 558598 -408
rect 558654 -464 558722 -408
rect 558778 -464 558846 -408
rect 558902 -464 589194 -408
rect 589250 -464 589318 -408
rect 589374 -464 589442 -408
rect 589498 -464 589566 -408
rect 589622 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect -956 -532 597020 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 5514 -532
rect 5570 -588 5638 -532
rect 5694 -588 5762 -532
rect 5818 -588 5886 -532
rect 5942 -588 36234 -532
rect 36290 -588 36358 -532
rect 36414 -588 36482 -532
rect 36538 -588 36606 -532
rect 36662 -588 66954 -532
rect 67010 -588 67078 -532
rect 67134 -588 67202 -532
rect 67258 -588 67326 -532
rect 67382 -588 97674 -532
rect 97730 -588 97798 -532
rect 97854 -588 97922 -532
rect 97978 -588 98046 -532
rect 98102 -588 128394 -532
rect 128450 -588 128518 -532
rect 128574 -588 128642 -532
rect 128698 -588 128766 -532
rect 128822 -588 159114 -532
rect 159170 -588 159238 -532
rect 159294 -588 159362 -532
rect 159418 -588 159486 -532
rect 159542 -588 189834 -532
rect 189890 -588 189958 -532
rect 190014 -588 190082 -532
rect 190138 -588 190206 -532
rect 190262 -588 220554 -532
rect 220610 -588 220678 -532
rect 220734 -588 220802 -532
rect 220858 -588 220926 -532
rect 220982 -588 251274 -532
rect 251330 -588 251398 -532
rect 251454 -588 251522 -532
rect 251578 -588 251646 -532
rect 251702 -588 281994 -532
rect 282050 -588 282118 -532
rect 282174 -588 282242 -532
rect 282298 -588 282366 -532
rect 282422 -588 312714 -532
rect 312770 -588 312838 -532
rect 312894 -588 312962 -532
rect 313018 -588 313086 -532
rect 313142 -588 343434 -532
rect 343490 -588 343558 -532
rect 343614 -588 343682 -532
rect 343738 -588 343806 -532
rect 343862 -588 374154 -532
rect 374210 -588 374278 -532
rect 374334 -588 374402 -532
rect 374458 -588 374526 -532
rect 374582 -588 404874 -532
rect 404930 -588 404998 -532
rect 405054 -588 405122 -532
rect 405178 -588 405246 -532
rect 405302 -588 435594 -532
rect 435650 -588 435718 -532
rect 435774 -588 435842 -532
rect 435898 -588 435966 -532
rect 436022 -588 466314 -532
rect 466370 -588 466438 -532
rect 466494 -588 466562 -532
rect 466618 -588 466686 -532
rect 466742 -588 497034 -532
rect 497090 -588 497158 -532
rect 497214 -588 497282 -532
rect 497338 -588 497406 -532
rect 497462 -588 527754 -532
rect 527810 -588 527878 -532
rect 527934 -588 528002 -532
rect 528058 -588 528126 -532
rect 528182 -588 558474 -532
rect 558530 -588 558598 -532
rect 558654 -588 558722 -532
rect 558778 -588 558846 -532
rect 558902 -588 589194 -532
rect 589250 -588 589318 -532
rect 589374 -588 589442 -532
rect 589498 -588 589566 -532
rect 589622 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect -956 -684 597020 -588
rect -1916 -1120 597980 -1024
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 592914 -1120
rect 592970 -1176 593038 -1120
rect 593094 -1176 593162 -1120
rect 593218 -1176 593286 -1120
rect 593342 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect -1916 -1244 597980 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 592914 -1244
rect 592970 -1300 593038 -1244
rect 593094 -1300 593162 -1244
rect 593218 -1300 593286 -1244
rect 593342 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect -1916 -1368 597980 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 592914 -1368
rect 592970 -1424 593038 -1368
rect 593094 -1424 593162 -1368
rect 593218 -1424 593286 -1368
rect 593342 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect -1916 -1492 597980 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 592914 -1492
rect 592970 -1548 593038 -1492
rect 593094 -1548 593162 -1492
rect 593218 -1548 593286 -1492
rect 593342 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect -1916 -1644 597980 -1548
use rift2Wrap  i_Rift2Wrap
timestamp 0
transform 1 0 8000 0 1 8000
box 0 0 574094 577678
<< labels >>
flabel metal3 s 595560 7112 597000 7336 0 FreeSans 896 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 595560 403592 597000 403816 0 FreeSans 896 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 595560 443240 597000 443464 0 FreeSans 896 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 595560 482888 597000 483112 0 FreeSans 896 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 595560 522536 597000 522760 0 FreeSans 896 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 595560 562184 597000 562408 0 FreeSans 896 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 584696 595560 584920 597000 0 FreeSans 896 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 518504 595560 518728 597000 0 FreeSans 896 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 452312 595560 452536 597000 0 FreeSans 896 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 386120 595560 386344 597000 0 FreeSans 896 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 319928 595560 320152 597000 0 FreeSans 896 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 595560 46760 597000 46984 0 FreeSans 896 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 253736 595560 253960 597000 0 FreeSans 896 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 187544 595560 187768 597000 0 FreeSans 896 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 121352 595560 121576 597000 0 FreeSans 896 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 55160 595560 55384 597000 0 FreeSans 896 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s -960 587160 480 587384 0 FreeSans 896 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s -960 544824 480 545048 0 FreeSans 896 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s -960 502488 480 502712 0 FreeSans 896 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s -960 460152 480 460376 0 FreeSans 896 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s -960 417816 480 418040 0 FreeSans 896 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s -960 375480 480 375704 0 FreeSans 896 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 595560 86408 597000 86632 0 FreeSans 896 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s -960 333144 480 333368 0 FreeSans 896 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s -960 290808 480 291032 0 FreeSans 896 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s -960 248472 480 248696 0 FreeSans 896 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s -960 206136 480 206360 0 FreeSans 896 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s -960 163800 480 164024 0 FreeSans 896 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s -960 121464 480 121688 0 FreeSans 896 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s -960 79128 480 79352 0 FreeSans 896 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s -960 36792 480 37016 0 FreeSans 896 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 595560 126056 597000 126280 0 FreeSans 896 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 595560 165704 597000 165928 0 FreeSans 896 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 595560 205352 597000 205576 0 FreeSans 896 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 595560 245000 597000 245224 0 FreeSans 896 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 595560 284648 597000 284872 0 FreeSans 896 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 595560 324296 597000 324520 0 FreeSans 896 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 595560 363944 597000 364168 0 FreeSans 896 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 595560 33544 597000 33768 0 FreeSans 896 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 595560 430024 597000 430248 0 FreeSans 896 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 595560 469672 597000 469896 0 FreeSans 896 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 595560 509320 597000 509544 0 FreeSans 896 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 595560 548968 597000 549192 0 FreeSans 896 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 595560 588616 597000 588840 0 FreeSans 896 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 540568 595560 540792 597000 0 FreeSans 896 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 474376 595560 474600 597000 0 FreeSans 896 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 408184 595560 408408 597000 0 FreeSans 896 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 341992 595560 342216 597000 0 FreeSans 896 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 275800 595560 276024 597000 0 FreeSans 896 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 595560 73192 597000 73416 0 FreeSans 896 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 209608 595560 209832 597000 0 FreeSans 896 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 143416 595560 143640 597000 0 FreeSans 896 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 77224 595560 77448 597000 0 FreeSans 896 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 11032 595560 11256 597000 0 FreeSans 896 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s -960 558936 480 559160 0 FreeSans 896 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s -960 516600 480 516824 0 FreeSans 896 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s -960 474264 480 474488 0 FreeSans 896 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s -960 431928 480 432152 0 FreeSans 896 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s -960 389592 480 389816 0 FreeSans 896 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s -960 347256 480 347480 0 FreeSans 896 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 595560 112840 597000 113064 0 FreeSans 896 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s -960 304920 480 305144 0 FreeSans 896 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s -960 262584 480 262808 0 FreeSans 896 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s -960 220248 480 220472 0 FreeSans 896 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s -960 177912 480 178136 0 FreeSans 896 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s -960 135576 480 135800 0 FreeSans 896 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s -960 93240 480 93464 0 FreeSans 896 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s -960 50904 480 51128 0 FreeSans 896 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s -960 8568 480 8792 0 FreeSans 896 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 595560 152488 597000 152712 0 FreeSans 896 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 595560 192136 597000 192360 0 FreeSans 896 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 595560 231784 597000 232008 0 FreeSans 896 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 595560 271432 597000 271656 0 FreeSans 896 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 595560 311080 597000 311304 0 FreeSans 896 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 595560 350728 597000 350952 0 FreeSans 896 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 595560 390376 597000 390600 0 FreeSans 896 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 595560 20328 597000 20552 0 FreeSans 896 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 595560 416808 597000 417032 0 FreeSans 896 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 595560 456456 597000 456680 0 FreeSans 896 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 595560 496104 597000 496328 0 FreeSans 896 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 595560 535752 597000 535976 0 FreeSans 896 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 595560 575400 597000 575624 0 FreeSans 896 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 562632 595560 562856 597000 0 FreeSans 896 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 496440 595560 496664 597000 0 FreeSans 896 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 430248 595560 430472 597000 0 FreeSans 896 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 364056 595560 364280 597000 0 FreeSans 896 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 297864 595560 298088 597000 0 FreeSans 896 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 595560 59976 597000 60200 0 FreeSans 896 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 231672 595560 231896 597000 0 FreeSans 896 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 165480 595560 165704 597000 0 FreeSans 896 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 99288 595560 99512 597000 0 FreeSans 896 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 33096 595560 33320 597000 0 FreeSans 896 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s -960 573048 480 573272 0 FreeSans 896 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s -960 530712 480 530936 0 FreeSans 896 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s -960 488376 480 488600 0 FreeSans 896 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s -960 446040 480 446264 0 FreeSans 896 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s -960 403704 480 403928 0 FreeSans 896 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s -960 361368 480 361592 0 FreeSans 896 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 595560 99624 597000 99848 0 FreeSans 896 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s -960 319032 480 319256 0 FreeSans 896 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s -960 276696 480 276920 0 FreeSans 896 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s -960 234360 480 234584 0 FreeSans 896 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s -960 192024 480 192248 0 FreeSans 896 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s -960 149688 480 149912 0 FreeSans 896 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s -960 107352 480 107576 0 FreeSans 896 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s -960 65016 480 65240 0 FreeSans 896 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s -960 22680 480 22904 0 FreeSans 896 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 595560 139272 597000 139496 0 FreeSans 896 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 595560 178920 597000 179144 0 FreeSans 896 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 595560 218568 597000 218792 0 FreeSans 896 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 595560 258216 597000 258440 0 FreeSans 896 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 595560 297864 597000 298088 0 FreeSans 896 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 595560 337512 597000 337736 0 FreeSans 896 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 595560 377160 597000 377384 0 FreeSans 896 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 213192 -960 213416 480 0 FreeSans 896 90 0 0 la_data_in[0]
port 114 nsew signal input
flabel metal2 s 270312 -960 270536 480 0 FreeSans 896 90 0 0 la_data_in[10]
port 115 nsew signal input
flabel metal2 s 276024 -960 276248 480 0 FreeSans 896 90 0 0 la_data_in[11]
port 116 nsew signal input
flabel metal2 s 281736 -960 281960 480 0 FreeSans 896 90 0 0 la_data_in[12]
port 117 nsew signal input
flabel metal2 s 287448 -960 287672 480 0 FreeSans 896 90 0 0 la_data_in[13]
port 118 nsew signal input
flabel metal2 s 293160 -960 293384 480 0 FreeSans 896 90 0 0 la_data_in[14]
port 119 nsew signal input
flabel metal2 s 298872 -960 299096 480 0 FreeSans 896 90 0 0 la_data_in[15]
port 120 nsew signal input
flabel metal2 s 304584 -960 304808 480 0 FreeSans 896 90 0 0 la_data_in[16]
port 121 nsew signal input
flabel metal2 s 310296 -960 310520 480 0 FreeSans 896 90 0 0 la_data_in[17]
port 122 nsew signal input
flabel metal2 s 316008 -960 316232 480 0 FreeSans 896 90 0 0 la_data_in[18]
port 123 nsew signal input
flabel metal2 s 321720 -960 321944 480 0 FreeSans 896 90 0 0 la_data_in[19]
port 124 nsew signal input
flabel metal2 s 218904 -960 219128 480 0 FreeSans 896 90 0 0 la_data_in[1]
port 125 nsew signal input
flabel metal2 s 327432 -960 327656 480 0 FreeSans 896 90 0 0 la_data_in[20]
port 126 nsew signal input
flabel metal2 s 333144 -960 333368 480 0 FreeSans 896 90 0 0 la_data_in[21]
port 127 nsew signal input
flabel metal2 s 338856 -960 339080 480 0 FreeSans 896 90 0 0 la_data_in[22]
port 128 nsew signal input
flabel metal2 s 344568 -960 344792 480 0 FreeSans 896 90 0 0 la_data_in[23]
port 129 nsew signal input
flabel metal2 s 350280 -960 350504 480 0 FreeSans 896 90 0 0 la_data_in[24]
port 130 nsew signal input
flabel metal2 s 355992 -960 356216 480 0 FreeSans 896 90 0 0 la_data_in[25]
port 131 nsew signal input
flabel metal2 s 361704 -960 361928 480 0 FreeSans 896 90 0 0 la_data_in[26]
port 132 nsew signal input
flabel metal2 s 367416 -960 367640 480 0 FreeSans 896 90 0 0 la_data_in[27]
port 133 nsew signal input
flabel metal2 s 373128 -960 373352 480 0 FreeSans 896 90 0 0 la_data_in[28]
port 134 nsew signal input
flabel metal2 s 378840 -960 379064 480 0 FreeSans 896 90 0 0 la_data_in[29]
port 135 nsew signal input
flabel metal2 s 224616 -960 224840 480 0 FreeSans 896 90 0 0 la_data_in[2]
port 136 nsew signal input
flabel metal2 s 384552 -960 384776 480 0 FreeSans 896 90 0 0 la_data_in[30]
port 137 nsew signal input
flabel metal2 s 390264 -960 390488 480 0 FreeSans 896 90 0 0 la_data_in[31]
port 138 nsew signal input
flabel metal2 s 395976 -960 396200 480 0 FreeSans 896 90 0 0 la_data_in[32]
port 139 nsew signal input
flabel metal2 s 401688 -960 401912 480 0 FreeSans 896 90 0 0 la_data_in[33]
port 140 nsew signal input
flabel metal2 s 407400 -960 407624 480 0 FreeSans 896 90 0 0 la_data_in[34]
port 141 nsew signal input
flabel metal2 s 413112 -960 413336 480 0 FreeSans 896 90 0 0 la_data_in[35]
port 142 nsew signal input
flabel metal2 s 418824 -960 419048 480 0 FreeSans 896 90 0 0 la_data_in[36]
port 143 nsew signal input
flabel metal2 s 424536 -960 424760 480 0 FreeSans 896 90 0 0 la_data_in[37]
port 144 nsew signal input
flabel metal2 s 430248 -960 430472 480 0 FreeSans 896 90 0 0 la_data_in[38]
port 145 nsew signal input
flabel metal2 s 435960 -960 436184 480 0 FreeSans 896 90 0 0 la_data_in[39]
port 146 nsew signal input
flabel metal2 s 230328 -960 230552 480 0 FreeSans 896 90 0 0 la_data_in[3]
port 147 nsew signal input
flabel metal2 s 441672 -960 441896 480 0 FreeSans 896 90 0 0 la_data_in[40]
port 148 nsew signal input
flabel metal2 s 447384 -960 447608 480 0 FreeSans 896 90 0 0 la_data_in[41]
port 149 nsew signal input
flabel metal2 s 453096 -960 453320 480 0 FreeSans 896 90 0 0 la_data_in[42]
port 150 nsew signal input
flabel metal2 s 458808 -960 459032 480 0 FreeSans 896 90 0 0 la_data_in[43]
port 151 nsew signal input
flabel metal2 s 464520 -960 464744 480 0 FreeSans 896 90 0 0 la_data_in[44]
port 152 nsew signal input
flabel metal2 s 470232 -960 470456 480 0 FreeSans 896 90 0 0 la_data_in[45]
port 153 nsew signal input
flabel metal2 s 475944 -960 476168 480 0 FreeSans 896 90 0 0 la_data_in[46]
port 154 nsew signal input
flabel metal2 s 481656 -960 481880 480 0 FreeSans 896 90 0 0 la_data_in[47]
port 155 nsew signal input
flabel metal2 s 487368 -960 487592 480 0 FreeSans 896 90 0 0 la_data_in[48]
port 156 nsew signal input
flabel metal2 s 493080 -960 493304 480 0 FreeSans 896 90 0 0 la_data_in[49]
port 157 nsew signal input
flabel metal2 s 236040 -960 236264 480 0 FreeSans 896 90 0 0 la_data_in[4]
port 158 nsew signal input
flabel metal2 s 498792 -960 499016 480 0 FreeSans 896 90 0 0 la_data_in[50]
port 159 nsew signal input
flabel metal2 s 504504 -960 504728 480 0 FreeSans 896 90 0 0 la_data_in[51]
port 160 nsew signal input
flabel metal2 s 510216 -960 510440 480 0 FreeSans 896 90 0 0 la_data_in[52]
port 161 nsew signal input
flabel metal2 s 515928 -960 516152 480 0 FreeSans 896 90 0 0 la_data_in[53]
port 162 nsew signal input
flabel metal2 s 521640 -960 521864 480 0 FreeSans 896 90 0 0 la_data_in[54]
port 163 nsew signal input
flabel metal2 s 527352 -960 527576 480 0 FreeSans 896 90 0 0 la_data_in[55]
port 164 nsew signal input
flabel metal2 s 533064 -960 533288 480 0 FreeSans 896 90 0 0 la_data_in[56]
port 165 nsew signal input
flabel metal2 s 538776 -960 539000 480 0 FreeSans 896 90 0 0 la_data_in[57]
port 166 nsew signal input
flabel metal2 s 544488 -960 544712 480 0 FreeSans 896 90 0 0 la_data_in[58]
port 167 nsew signal input
flabel metal2 s 550200 -960 550424 480 0 FreeSans 896 90 0 0 la_data_in[59]
port 168 nsew signal input
flabel metal2 s 241752 -960 241976 480 0 FreeSans 896 90 0 0 la_data_in[5]
port 169 nsew signal input
flabel metal2 s 555912 -960 556136 480 0 FreeSans 896 90 0 0 la_data_in[60]
port 170 nsew signal input
flabel metal2 s 561624 -960 561848 480 0 FreeSans 896 90 0 0 la_data_in[61]
port 171 nsew signal input
flabel metal2 s 567336 -960 567560 480 0 FreeSans 896 90 0 0 la_data_in[62]
port 172 nsew signal input
flabel metal2 s 573048 -960 573272 480 0 FreeSans 896 90 0 0 la_data_in[63]
port 173 nsew signal input
flabel metal2 s 247464 -960 247688 480 0 FreeSans 896 90 0 0 la_data_in[6]
port 174 nsew signal input
flabel metal2 s 253176 -960 253400 480 0 FreeSans 896 90 0 0 la_data_in[7]
port 175 nsew signal input
flabel metal2 s 258888 -960 259112 480 0 FreeSans 896 90 0 0 la_data_in[8]
port 176 nsew signal input
flabel metal2 s 264600 -960 264824 480 0 FreeSans 896 90 0 0 la_data_in[9]
port 177 nsew signal input
flabel metal2 s 215096 -960 215320 480 0 FreeSans 896 90 0 0 la_data_out[0]
port 178 nsew signal tristate
flabel metal2 s 272216 -960 272440 480 0 FreeSans 896 90 0 0 la_data_out[10]
port 179 nsew signal tristate
flabel metal2 s 277928 -960 278152 480 0 FreeSans 896 90 0 0 la_data_out[11]
port 180 nsew signal tristate
flabel metal2 s 283640 -960 283864 480 0 FreeSans 896 90 0 0 la_data_out[12]
port 181 nsew signal tristate
flabel metal2 s 289352 -960 289576 480 0 FreeSans 896 90 0 0 la_data_out[13]
port 182 nsew signal tristate
flabel metal2 s 295064 -960 295288 480 0 FreeSans 896 90 0 0 la_data_out[14]
port 183 nsew signal tristate
flabel metal2 s 300776 -960 301000 480 0 FreeSans 896 90 0 0 la_data_out[15]
port 184 nsew signal tristate
flabel metal2 s 306488 -960 306712 480 0 FreeSans 896 90 0 0 la_data_out[16]
port 185 nsew signal tristate
flabel metal2 s 312200 -960 312424 480 0 FreeSans 896 90 0 0 la_data_out[17]
port 186 nsew signal tristate
flabel metal2 s 317912 -960 318136 480 0 FreeSans 896 90 0 0 la_data_out[18]
port 187 nsew signal tristate
flabel metal2 s 323624 -960 323848 480 0 FreeSans 896 90 0 0 la_data_out[19]
port 188 nsew signal tristate
flabel metal2 s 220808 -960 221032 480 0 FreeSans 896 90 0 0 la_data_out[1]
port 189 nsew signal tristate
flabel metal2 s 329336 -960 329560 480 0 FreeSans 896 90 0 0 la_data_out[20]
port 190 nsew signal tristate
flabel metal2 s 335048 -960 335272 480 0 FreeSans 896 90 0 0 la_data_out[21]
port 191 nsew signal tristate
flabel metal2 s 340760 -960 340984 480 0 FreeSans 896 90 0 0 la_data_out[22]
port 192 nsew signal tristate
flabel metal2 s 346472 -960 346696 480 0 FreeSans 896 90 0 0 la_data_out[23]
port 193 nsew signal tristate
flabel metal2 s 352184 -960 352408 480 0 FreeSans 896 90 0 0 la_data_out[24]
port 194 nsew signal tristate
flabel metal2 s 357896 -960 358120 480 0 FreeSans 896 90 0 0 la_data_out[25]
port 195 nsew signal tristate
flabel metal2 s 363608 -960 363832 480 0 FreeSans 896 90 0 0 la_data_out[26]
port 196 nsew signal tristate
flabel metal2 s 369320 -960 369544 480 0 FreeSans 896 90 0 0 la_data_out[27]
port 197 nsew signal tristate
flabel metal2 s 375032 -960 375256 480 0 FreeSans 896 90 0 0 la_data_out[28]
port 198 nsew signal tristate
flabel metal2 s 380744 -960 380968 480 0 FreeSans 896 90 0 0 la_data_out[29]
port 199 nsew signal tristate
flabel metal2 s 226520 -960 226744 480 0 FreeSans 896 90 0 0 la_data_out[2]
port 200 nsew signal tristate
flabel metal2 s 386456 -960 386680 480 0 FreeSans 896 90 0 0 la_data_out[30]
port 201 nsew signal tristate
flabel metal2 s 392168 -960 392392 480 0 FreeSans 896 90 0 0 la_data_out[31]
port 202 nsew signal tristate
flabel metal2 s 397880 -960 398104 480 0 FreeSans 896 90 0 0 la_data_out[32]
port 203 nsew signal tristate
flabel metal2 s 403592 -960 403816 480 0 FreeSans 896 90 0 0 la_data_out[33]
port 204 nsew signal tristate
flabel metal2 s 409304 -960 409528 480 0 FreeSans 896 90 0 0 la_data_out[34]
port 205 nsew signal tristate
flabel metal2 s 415016 -960 415240 480 0 FreeSans 896 90 0 0 la_data_out[35]
port 206 nsew signal tristate
flabel metal2 s 420728 -960 420952 480 0 FreeSans 896 90 0 0 la_data_out[36]
port 207 nsew signal tristate
flabel metal2 s 426440 -960 426664 480 0 FreeSans 896 90 0 0 la_data_out[37]
port 208 nsew signal tristate
flabel metal2 s 432152 -960 432376 480 0 FreeSans 896 90 0 0 la_data_out[38]
port 209 nsew signal tristate
flabel metal2 s 437864 -960 438088 480 0 FreeSans 896 90 0 0 la_data_out[39]
port 210 nsew signal tristate
flabel metal2 s 232232 -960 232456 480 0 FreeSans 896 90 0 0 la_data_out[3]
port 211 nsew signal tristate
flabel metal2 s 443576 -960 443800 480 0 FreeSans 896 90 0 0 la_data_out[40]
port 212 nsew signal tristate
flabel metal2 s 449288 -960 449512 480 0 FreeSans 896 90 0 0 la_data_out[41]
port 213 nsew signal tristate
flabel metal2 s 455000 -960 455224 480 0 FreeSans 896 90 0 0 la_data_out[42]
port 214 nsew signal tristate
flabel metal2 s 460712 -960 460936 480 0 FreeSans 896 90 0 0 la_data_out[43]
port 215 nsew signal tristate
flabel metal2 s 466424 -960 466648 480 0 FreeSans 896 90 0 0 la_data_out[44]
port 216 nsew signal tristate
flabel metal2 s 472136 -960 472360 480 0 FreeSans 896 90 0 0 la_data_out[45]
port 217 nsew signal tristate
flabel metal2 s 477848 -960 478072 480 0 FreeSans 896 90 0 0 la_data_out[46]
port 218 nsew signal tristate
flabel metal2 s 483560 -960 483784 480 0 FreeSans 896 90 0 0 la_data_out[47]
port 219 nsew signal tristate
flabel metal2 s 489272 -960 489496 480 0 FreeSans 896 90 0 0 la_data_out[48]
port 220 nsew signal tristate
flabel metal2 s 494984 -960 495208 480 0 FreeSans 896 90 0 0 la_data_out[49]
port 221 nsew signal tristate
flabel metal2 s 237944 -960 238168 480 0 FreeSans 896 90 0 0 la_data_out[4]
port 222 nsew signal tristate
flabel metal2 s 500696 -960 500920 480 0 FreeSans 896 90 0 0 la_data_out[50]
port 223 nsew signal tristate
flabel metal2 s 506408 -960 506632 480 0 FreeSans 896 90 0 0 la_data_out[51]
port 224 nsew signal tristate
flabel metal2 s 512120 -960 512344 480 0 FreeSans 896 90 0 0 la_data_out[52]
port 225 nsew signal tristate
flabel metal2 s 517832 -960 518056 480 0 FreeSans 896 90 0 0 la_data_out[53]
port 226 nsew signal tristate
flabel metal2 s 523544 -960 523768 480 0 FreeSans 896 90 0 0 la_data_out[54]
port 227 nsew signal tristate
flabel metal2 s 529256 -960 529480 480 0 FreeSans 896 90 0 0 la_data_out[55]
port 228 nsew signal tristate
flabel metal2 s 534968 -960 535192 480 0 FreeSans 896 90 0 0 la_data_out[56]
port 229 nsew signal tristate
flabel metal2 s 540680 -960 540904 480 0 FreeSans 896 90 0 0 la_data_out[57]
port 230 nsew signal tristate
flabel metal2 s 546392 -960 546616 480 0 FreeSans 896 90 0 0 la_data_out[58]
port 231 nsew signal tristate
flabel metal2 s 552104 -960 552328 480 0 FreeSans 896 90 0 0 la_data_out[59]
port 232 nsew signal tristate
flabel metal2 s 243656 -960 243880 480 0 FreeSans 896 90 0 0 la_data_out[5]
port 233 nsew signal tristate
flabel metal2 s 557816 -960 558040 480 0 FreeSans 896 90 0 0 la_data_out[60]
port 234 nsew signal tristate
flabel metal2 s 563528 -960 563752 480 0 FreeSans 896 90 0 0 la_data_out[61]
port 235 nsew signal tristate
flabel metal2 s 569240 -960 569464 480 0 FreeSans 896 90 0 0 la_data_out[62]
port 236 nsew signal tristate
flabel metal2 s 574952 -960 575176 480 0 FreeSans 896 90 0 0 la_data_out[63]
port 237 nsew signal tristate
flabel metal2 s 249368 -960 249592 480 0 FreeSans 896 90 0 0 la_data_out[6]
port 238 nsew signal tristate
flabel metal2 s 255080 -960 255304 480 0 FreeSans 896 90 0 0 la_data_out[7]
port 239 nsew signal tristate
flabel metal2 s 260792 -960 261016 480 0 FreeSans 896 90 0 0 la_data_out[8]
port 240 nsew signal tristate
flabel metal2 s 266504 -960 266728 480 0 FreeSans 896 90 0 0 la_data_out[9]
port 241 nsew signal tristate
flabel metal2 s 217000 -960 217224 480 0 FreeSans 896 90 0 0 la_oenb[0]
port 242 nsew signal input
flabel metal2 s 274120 -960 274344 480 0 FreeSans 896 90 0 0 la_oenb[10]
port 243 nsew signal input
flabel metal2 s 279832 -960 280056 480 0 FreeSans 896 90 0 0 la_oenb[11]
port 244 nsew signal input
flabel metal2 s 285544 -960 285768 480 0 FreeSans 896 90 0 0 la_oenb[12]
port 245 nsew signal input
flabel metal2 s 291256 -960 291480 480 0 FreeSans 896 90 0 0 la_oenb[13]
port 246 nsew signal input
flabel metal2 s 296968 -960 297192 480 0 FreeSans 896 90 0 0 la_oenb[14]
port 247 nsew signal input
flabel metal2 s 302680 -960 302904 480 0 FreeSans 896 90 0 0 la_oenb[15]
port 248 nsew signal input
flabel metal2 s 308392 -960 308616 480 0 FreeSans 896 90 0 0 la_oenb[16]
port 249 nsew signal input
flabel metal2 s 314104 -960 314328 480 0 FreeSans 896 90 0 0 la_oenb[17]
port 250 nsew signal input
flabel metal2 s 319816 -960 320040 480 0 FreeSans 896 90 0 0 la_oenb[18]
port 251 nsew signal input
flabel metal2 s 325528 -960 325752 480 0 FreeSans 896 90 0 0 la_oenb[19]
port 252 nsew signal input
flabel metal2 s 222712 -960 222936 480 0 FreeSans 896 90 0 0 la_oenb[1]
port 253 nsew signal input
flabel metal2 s 331240 -960 331464 480 0 FreeSans 896 90 0 0 la_oenb[20]
port 254 nsew signal input
flabel metal2 s 336952 -960 337176 480 0 FreeSans 896 90 0 0 la_oenb[21]
port 255 nsew signal input
flabel metal2 s 342664 -960 342888 480 0 FreeSans 896 90 0 0 la_oenb[22]
port 256 nsew signal input
flabel metal2 s 348376 -960 348600 480 0 FreeSans 896 90 0 0 la_oenb[23]
port 257 nsew signal input
flabel metal2 s 354088 -960 354312 480 0 FreeSans 896 90 0 0 la_oenb[24]
port 258 nsew signal input
flabel metal2 s 359800 -960 360024 480 0 FreeSans 896 90 0 0 la_oenb[25]
port 259 nsew signal input
flabel metal2 s 365512 -960 365736 480 0 FreeSans 896 90 0 0 la_oenb[26]
port 260 nsew signal input
flabel metal2 s 371224 -960 371448 480 0 FreeSans 896 90 0 0 la_oenb[27]
port 261 nsew signal input
flabel metal2 s 376936 -960 377160 480 0 FreeSans 896 90 0 0 la_oenb[28]
port 262 nsew signal input
flabel metal2 s 382648 -960 382872 480 0 FreeSans 896 90 0 0 la_oenb[29]
port 263 nsew signal input
flabel metal2 s 228424 -960 228648 480 0 FreeSans 896 90 0 0 la_oenb[2]
port 264 nsew signal input
flabel metal2 s 388360 -960 388584 480 0 FreeSans 896 90 0 0 la_oenb[30]
port 265 nsew signal input
flabel metal2 s 394072 -960 394296 480 0 FreeSans 896 90 0 0 la_oenb[31]
port 266 nsew signal input
flabel metal2 s 399784 -960 400008 480 0 FreeSans 896 90 0 0 la_oenb[32]
port 267 nsew signal input
flabel metal2 s 405496 -960 405720 480 0 FreeSans 896 90 0 0 la_oenb[33]
port 268 nsew signal input
flabel metal2 s 411208 -960 411432 480 0 FreeSans 896 90 0 0 la_oenb[34]
port 269 nsew signal input
flabel metal2 s 416920 -960 417144 480 0 FreeSans 896 90 0 0 la_oenb[35]
port 270 nsew signal input
flabel metal2 s 422632 -960 422856 480 0 FreeSans 896 90 0 0 la_oenb[36]
port 271 nsew signal input
flabel metal2 s 428344 -960 428568 480 0 FreeSans 896 90 0 0 la_oenb[37]
port 272 nsew signal input
flabel metal2 s 434056 -960 434280 480 0 FreeSans 896 90 0 0 la_oenb[38]
port 273 nsew signal input
flabel metal2 s 439768 -960 439992 480 0 FreeSans 896 90 0 0 la_oenb[39]
port 274 nsew signal input
flabel metal2 s 234136 -960 234360 480 0 FreeSans 896 90 0 0 la_oenb[3]
port 275 nsew signal input
flabel metal2 s 445480 -960 445704 480 0 FreeSans 896 90 0 0 la_oenb[40]
port 276 nsew signal input
flabel metal2 s 451192 -960 451416 480 0 FreeSans 896 90 0 0 la_oenb[41]
port 277 nsew signal input
flabel metal2 s 456904 -960 457128 480 0 FreeSans 896 90 0 0 la_oenb[42]
port 278 nsew signal input
flabel metal2 s 462616 -960 462840 480 0 FreeSans 896 90 0 0 la_oenb[43]
port 279 nsew signal input
flabel metal2 s 468328 -960 468552 480 0 FreeSans 896 90 0 0 la_oenb[44]
port 280 nsew signal input
flabel metal2 s 474040 -960 474264 480 0 FreeSans 896 90 0 0 la_oenb[45]
port 281 nsew signal input
flabel metal2 s 479752 -960 479976 480 0 FreeSans 896 90 0 0 la_oenb[46]
port 282 nsew signal input
flabel metal2 s 485464 -960 485688 480 0 FreeSans 896 90 0 0 la_oenb[47]
port 283 nsew signal input
flabel metal2 s 491176 -960 491400 480 0 FreeSans 896 90 0 0 la_oenb[48]
port 284 nsew signal input
flabel metal2 s 496888 -960 497112 480 0 FreeSans 896 90 0 0 la_oenb[49]
port 285 nsew signal input
flabel metal2 s 239848 -960 240072 480 0 FreeSans 896 90 0 0 la_oenb[4]
port 286 nsew signal input
flabel metal2 s 502600 -960 502824 480 0 FreeSans 896 90 0 0 la_oenb[50]
port 287 nsew signal input
flabel metal2 s 508312 -960 508536 480 0 FreeSans 896 90 0 0 la_oenb[51]
port 288 nsew signal input
flabel metal2 s 514024 -960 514248 480 0 FreeSans 896 90 0 0 la_oenb[52]
port 289 nsew signal input
flabel metal2 s 519736 -960 519960 480 0 FreeSans 896 90 0 0 la_oenb[53]
port 290 nsew signal input
flabel metal2 s 525448 -960 525672 480 0 FreeSans 896 90 0 0 la_oenb[54]
port 291 nsew signal input
flabel metal2 s 531160 -960 531384 480 0 FreeSans 896 90 0 0 la_oenb[55]
port 292 nsew signal input
flabel metal2 s 536872 -960 537096 480 0 FreeSans 896 90 0 0 la_oenb[56]
port 293 nsew signal input
flabel metal2 s 542584 -960 542808 480 0 FreeSans 896 90 0 0 la_oenb[57]
port 294 nsew signal input
flabel metal2 s 548296 -960 548520 480 0 FreeSans 896 90 0 0 la_oenb[58]
port 295 nsew signal input
flabel metal2 s 554008 -960 554232 480 0 FreeSans 896 90 0 0 la_oenb[59]
port 296 nsew signal input
flabel metal2 s 245560 -960 245784 480 0 FreeSans 896 90 0 0 la_oenb[5]
port 297 nsew signal input
flabel metal2 s 559720 -960 559944 480 0 FreeSans 896 90 0 0 la_oenb[60]
port 298 nsew signal input
flabel metal2 s 565432 -960 565656 480 0 FreeSans 896 90 0 0 la_oenb[61]
port 299 nsew signal input
flabel metal2 s 571144 -960 571368 480 0 FreeSans 896 90 0 0 la_oenb[62]
port 300 nsew signal input
flabel metal2 s 576856 -960 577080 480 0 FreeSans 896 90 0 0 la_oenb[63]
port 301 nsew signal input
flabel metal2 s 251272 -960 251496 480 0 FreeSans 896 90 0 0 la_oenb[6]
port 302 nsew signal input
flabel metal2 s 256984 -960 257208 480 0 FreeSans 896 90 0 0 la_oenb[7]
port 303 nsew signal input
flabel metal2 s 262696 -960 262920 480 0 FreeSans 896 90 0 0 la_oenb[8]
port 304 nsew signal input
flabel metal2 s 268408 -960 268632 480 0 FreeSans 896 90 0 0 la_oenb[9]
port 305 nsew signal input
flabel metal2 s 578760 -960 578984 480 0 FreeSans 896 90 0 0 user_clock2
port 306 nsew signal input
flabel metal2 s 580664 -960 580888 480 0 FreeSans 896 90 0 0 user_irq[0]
port 307 nsew signal tristate
flabel metal2 s 582568 -960 582792 480 0 FreeSans 896 90 0 0 user_irq[1]
port 308 nsew signal tristate
flabel metal2 s 584472 -960 584696 480 0 FreeSans 896 90 0 0 user_irq[2]
port 309 nsew signal tristate
flabel metal4 s -956 -684 -336 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 -684 597020 -64 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 596688 597020 597308 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 596400 -684 597020 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 5418 -1644 6038 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 36138 -1644 36758 7250 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 -1644 67478 7250 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 97578 -1644 98198 7250 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 128298 -1644 128918 7250 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 159018 -1644 159638 7250 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 189738 -1644 190358 7250 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 -1644 221078 7250 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 -1644 251798 7250 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 281898 -1644 282518 7250 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 -1644 313238 7250 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 343338 -1644 343958 7250 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 374058 -1644 374678 7250 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 404778 -1644 405398 7250 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435498 -1644 436118 7250 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 466218 -1644 466838 7250 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 496938 -1644 497558 7250 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 527658 -1644 528278 7250 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 558378 -1644 558998 7250 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 589098 -1644 589718 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 3826 597980 4446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 21826 597980 22446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 39826 597980 40446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 57826 597980 58446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 75826 597980 76446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 93826 597980 94446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 111826 597980 112446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 129826 597980 130446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 147826 597980 148446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 165826 597980 166446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 183826 597980 184446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 201826 597980 202446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 219826 597980 220446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 237826 597980 238446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 255826 597980 256446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 273826 597980 274446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 291826 597980 292446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 309826 597980 310446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 327826 597980 328446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 345826 597980 346446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 363826 597980 364446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 381826 597980 382446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 399826 597980 400446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 417826 597980 418446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 435826 597980 436446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 453826 597980 454446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 471826 597980 472446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 489826 597980 490446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 507826 597980 508446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 525826 597980 526446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 543826 597980 544446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 561826 597980 562446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 579826 597980 580446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s -1916 -1644 -1296 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 -1644 597980 -1024 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 597648 597980 598268 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 597360 -1644 597980 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 9138 584990 9758 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 39858 584990 40478 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 584990 71198 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 101298 584990 101918 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132018 584990 132638 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 584990 163358 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 193458 584990 194078 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 584990 224798 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 254898 584990 255518 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 285618 584990 286238 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 584990 316958 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 347058 584990 347678 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 377778 584990 378398 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 408498 584990 409118 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 439218 584990 439838 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 469938 584990 470558 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 500658 584990 501278 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 531378 584990 531998 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 562098 584990 562718 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 592818 -1644 593438 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 9826 597980 10446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 27826 597980 28446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 45826 597980 46446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 63826 597980 64446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 81826 597980 82446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 99826 597980 100446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 117826 597980 118446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 135826 597980 136446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 153826 597980 154446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 171826 597980 172446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 189826 597980 190446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 207826 597980 208446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 225826 597980 226446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 243826 597980 244446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 261826 597980 262446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 279826 597980 280446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 297826 597980 298446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 315826 597980 316446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 333826 597980 334446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 351826 597980 352446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 369826 597980 370446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 387826 597980 388446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 405826 597980 406446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 423826 597980 424446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 441826 597980 442446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 459826 597980 460446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 477826 597980 478446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 495826 597980 496446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 513826 597980 514446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 531826 597980 532446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 549826 597980 550446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 567826 597980 568446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 585826 597980 586446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal2 s 11368 -960 11592 480 0 FreeSans 896 90 0 0 wb_clk_i
port 312 nsew signal input
flabel metal2 s 13272 -960 13496 480 0 FreeSans 896 90 0 0 wb_rst_i
port 313 nsew signal input
flabel metal2 s 15176 -960 15400 480 0 FreeSans 896 90 0 0 wbs_ack_o
port 314 nsew signal tristate
flabel metal2 s 22792 -960 23016 480 0 FreeSans 896 90 0 0 wbs_adr_i[0]
port 315 nsew signal input
flabel metal2 s 87528 -960 87752 480 0 FreeSans 896 90 0 0 wbs_adr_i[10]
port 316 nsew signal input
flabel metal2 s 93240 -960 93464 480 0 FreeSans 896 90 0 0 wbs_adr_i[11]
port 317 nsew signal input
flabel metal2 s 98952 -960 99176 480 0 FreeSans 896 90 0 0 wbs_adr_i[12]
port 318 nsew signal input
flabel metal2 s 104664 -960 104888 480 0 FreeSans 896 90 0 0 wbs_adr_i[13]
port 319 nsew signal input
flabel metal2 s 110376 -960 110600 480 0 FreeSans 896 90 0 0 wbs_adr_i[14]
port 320 nsew signal input
flabel metal2 s 116088 -960 116312 480 0 FreeSans 896 90 0 0 wbs_adr_i[15]
port 321 nsew signal input
flabel metal2 s 121800 -960 122024 480 0 FreeSans 896 90 0 0 wbs_adr_i[16]
port 322 nsew signal input
flabel metal2 s 127512 -960 127736 480 0 FreeSans 896 90 0 0 wbs_adr_i[17]
port 323 nsew signal input
flabel metal2 s 133224 -960 133448 480 0 FreeSans 896 90 0 0 wbs_adr_i[18]
port 324 nsew signal input
flabel metal2 s 138936 -960 139160 480 0 FreeSans 896 90 0 0 wbs_adr_i[19]
port 325 nsew signal input
flabel metal2 s 30408 -960 30632 480 0 FreeSans 896 90 0 0 wbs_adr_i[1]
port 326 nsew signal input
flabel metal2 s 144648 -960 144872 480 0 FreeSans 896 90 0 0 wbs_adr_i[20]
port 327 nsew signal input
flabel metal2 s 150360 -960 150584 480 0 FreeSans 896 90 0 0 wbs_adr_i[21]
port 328 nsew signal input
flabel metal2 s 156072 -960 156296 480 0 FreeSans 896 90 0 0 wbs_adr_i[22]
port 329 nsew signal input
flabel metal2 s 161784 -960 162008 480 0 FreeSans 896 90 0 0 wbs_adr_i[23]
port 330 nsew signal input
flabel metal2 s 167496 -960 167720 480 0 FreeSans 896 90 0 0 wbs_adr_i[24]
port 331 nsew signal input
flabel metal2 s 173208 -960 173432 480 0 FreeSans 896 90 0 0 wbs_adr_i[25]
port 332 nsew signal input
flabel metal2 s 178920 -960 179144 480 0 FreeSans 896 90 0 0 wbs_adr_i[26]
port 333 nsew signal input
flabel metal2 s 184632 -960 184856 480 0 FreeSans 896 90 0 0 wbs_adr_i[27]
port 334 nsew signal input
flabel metal2 s 190344 -960 190568 480 0 FreeSans 896 90 0 0 wbs_adr_i[28]
port 335 nsew signal input
flabel metal2 s 196056 -960 196280 480 0 FreeSans 896 90 0 0 wbs_adr_i[29]
port 336 nsew signal input
flabel metal2 s 38024 -960 38248 480 0 FreeSans 896 90 0 0 wbs_adr_i[2]
port 337 nsew signal input
flabel metal2 s 201768 -960 201992 480 0 FreeSans 896 90 0 0 wbs_adr_i[30]
port 338 nsew signal input
flabel metal2 s 207480 -960 207704 480 0 FreeSans 896 90 0 0 wbs_adr_i[31]
port 339 nsew signal input
flabel metal2 s 45640 -960 45864 480 0 FreeSans 896 90 0 0 wbs_adr_i[3]
port 340 nsew signal input
flabel metal2 s 53256 -960 53480 480 0 FreeSans 896 90 0 0 wbs_adr_i[4]
port 341 nsew signal input
flabel metal2 s 58968 -960 59192 480 0 FreeSans 896 90 0 0 wbs_adr_i[5]
port 342 nsew signal input
flabel metal2 s 64680 -960 64904 480 0 FreeSans 896 90 0 0 wbs_adr_i[6]
port 343 nsew signal input
flabel metal2 s 70392 -960 70616 480 0 FreeSans 896 90 0 0 wbs_adr_i[7]
port 344 nsew signal input
flabel metal2 s 76104 -960 76328 480 0 FreeSans 896 90 0 0 wbs_adr_i[8]
port 345 nsew signal input
flabel metal2 s 81816 -960 82040 480 0 FreeSans 896 90 0 0 wbs_adr_i[9]
port 346 nsew signal input
flabel metal2 s 17080 -960 17304 480 0 FreeSans 896 90 0 0 wbs_cyc_i
port 347 nsew signal input
flabel metal2 s 24696 -960 24920 480 0 FreeSans 896 90 0 0 wbs_dat_i[0]
port 348 nsew signal input
flabel metal2 s 89432 -960 89656 480 0 FreeSans 896 90 0 0 wbs_dat_i[10]
port 349 nsew signal input
flabel metal2 s 95144 -960 95368 480 0 FreeSans 896 90 0 0 wbs_dat_i[11]
port 350 nsew signal input
flabel metal2 s 100856 -960 101080 480 0 FreeSans 896 90 0 0 wbs_dat_i[12]
port 351 nsew signal input
flabel metal2 s 106568 -960 106792 480 0 FreeSans 896 90 0 0 wbs_dat_i[13]
port 352 nsew signal input
flabel metal2 s 112280 -960 112504 480 0 FreeSans 896 90 0 0 wbs_dat_i[14]
port 353 nsew signal input
flabel metal2 s 117992 -960 118216 480 0 FreeSans 896 90 0 0 wbs_dat_i[15]
port 354 nsew signal input
flabel metal2 s 123704 -960 123928 480 0 FreeSans 896 90 0 0 wbs_dat_i[16]
port 355 nsew signal input
flabel metal2 s 129416 -960 129640 480 0 FreeSans 896 90 0 0 wbs_dat_i[17]
port 356 nsew signal input
flabel metal2 s 135128 -960 135352 480 0 FreeSans 896 90 0 0 wbs_dat_i[18]
port 357 nsew signal input
flabel metal2 s 140840 -960 141064 480 0 FreeSans 896 90 0 0 wbs_dat_i[19]
port 358 nsew signal input
flabel metal2 s 32312 -960 32536 480 0 FreeSans 896 90 0 0 wbs_dat_i[1]
port 359 nsew signal input
flabel metal2 s 146552 -960 146776 480 0 FreeSans 896 90 0 0 wbs_dat_i[20]
port 360 nsew signal input
flabel metal2 s 152264 -960 152488 480 0 FreeSans 896 90 0 0 wbs_dat_i[21]
port 361 nsew signal input
flabel metal2 s 157976 -960 158200 480 0 FreeSans 896 90 0 0 wbs_dat_i[22]
port 362 nsew signal input
flabel metal2 s 163688 -960 163912 480 0 FreeSans 896 90 0 0 wbs_dat_i[23]
port 363 nsew signal input
flabel metal2 s 169400 -960 169624 480 0 FreeSans 896 90 0 0 wbs_dat_i[24]
port 364 nsew signal input
flabel metal2 s 175112 -960 175336 480 0 FreeSans 896 90 0 0 wbs_dat_i[25]
port 365 nsew signal input
flabel metal2 s 180824 -960 181048 480 0 FreeSans 896 90 0 0 wbs_dat_i[26]
port 366 nsew signal input
flabel metal2 s 186536 -960 186760 480 0 FreeSans 896 90 0 0 wbs_dat_i[27]
port 367 nsew signal input
flabel metal2 s 192248 -960 192472 480 0 FreeSans 896 90 0 0 wbs_dat_i[28]
port 368 nsew signal input
flabel metal2 s 197960 -960 198184 480 0 FreeSans 896 90 0 0 wbs_dat_i[29]
port 369 nsew signal input
flabel metal2 s 39928 -960 40152 480 0 FreeSans 896 90 0 0 wbs_dat_i[2]
port 370 nsew signal input
flabel metal2 s 203672 -960 203896 480 0 FreeSans 896 90 0 0 wbs_dat_i[30]
port 371 nsew signal input
flabel metal2 s 209384 -960 209608 480 0 FreeSans 896 90 0 0 wbs_dat_i[31]
port 372 nsew signal input
flabel metal2 s 47544 -960 47768 480 0 FreeSans 896 90 0 0 wbs_dat_i[3]
port 373 nsew signal input
flabel metal2 s 55160 -960 55384 480 0 FreeSans 896 90 0 0 wbs_dat_i[4]
port 374 nsew signal input
flabel metal2 s 60872 -960 61096 480 0 FreeSans 896 90 0 0 wbs_dat_i[5]
port 375 nsew signal input
flabel metal2 s 66584 -960 66808 480 0 FreeSans 896 90 0 0 wbs_dat_i[6]
port 376 nsew signal input
flabel metal2 s 72296 -960 72520 480 0 FreeSans 896 90 0 0 wbs_dat_i[7]
port 377 nsew signal input
flabel metal2 s 78008 -960 78232 480 0 FreeSans 896 90 0 0 wbs_dat_i[8]
port 378 nsew signal input
flabel metal2 s 83720 -960 83944 480 0 FreeSans 896 90 0 0 wbs_dat_i[9]
port 379 nsew signal input
flabel metal2 s 26600 -960 26824 480 0 FreeSans 896 90 0 0 wbs_dat_o[0]
port 380 nsew signal tristate
flabel metal2 s 91336 -960 91560 480 0 FreeSans 896 90 0 0 wbs_dat_o[10]
port 381 nsew signal tristate
flabel metal2 s 97048 -960 97272 480 0 FreeSans 896 90 0 0 wbs_dat_o[11]
port 382 nsew signal tristate
flabel metal2 s 102760 -960 102984 480 0 FreeSans 896 90 0 0 wbs_dat_o[12]
port 383 nsew signal tristate
flabel metal2 s 108472 -960 108696 480 0 FreeSans 896 90 0 0 wbs_dat_o[13]
port 384 nsew signal tristate
flabel metal2 s 114184 -960 114408 480 0 FreeSans 896 90 0 0 wbs_dat_o[14]
port 385 nsew signal tristate
flabel metal2 s 119896 -960 120120 480 0 FreeSans 896 90 0 0 wbs_dat_o[15]
port 386 nsew signal tristate
flabel metal2 s 125608 -960 125832 480 0 FreeSans 896 90 0 0 wbs_dat_o[16]
port 387 nsew signal tristate
flabel metal2 s 131320 -960 131544 480 0 FreeSans 896 90 0 0 wbs_dat_o[17]
port 388 nsew signal tristate
flabel metal2 s 137032 -960 137256 480 0 FreeSans 896 90 0 0 wbs_dat_o[18]
port 389 nsew signal tristate
flabel metal2 s 142744 -960 142968 480 0 FreeSans 896 90 0 0 wbs_dat_o[19]
port 390 nsew signal tristate
flabel metal2 s 34216 -960 34440 480 0 FreeSans 896 90 0 0 wbs_dat_o[1]
port 391 nsew signal tristate
flabel metal2 s 148456 -960 148680 480 0 FreeSans 896 90 0 0 wbs_dat_o[20]
port 392 nsew signal tristate
flabel metal2 s 154168 -960 154392 480 0 FreeSans 896 90 0 0 wbs_dat_o[21]
port 393 nsew signal tristate
flabel metal2 s 159880 -960 160104 480 0 FreeSans 896 90 0 0 wbs_dat_o[22]
port 394 nsew signal tristate
flabel metal2 s 165592 -960 165816 480 0 FreeSans 896 90 0 0 wbs_dat_o[23]
port 395 nsew signal tristate
flabel metal2 s 171304 -960 171528 480 0 FreeSans 896 90 0 0 wbs_dat_o[24]
port 396 nsew signal tristate
flabel metal2 s 177016 -960 177240 480 0 FreeSans 896 90 0 0 wbs_dat_o[25]
port 397 nsew signal tristate
flabel metal2 s 182728 -960 182952 480 0 FreeSans 896 90 0 0 wbs_dat_o[26]
port 398 nsew signal tristate
flabel metal2 s 188440 -960 188664 480 0 FreeSans 896 90 0 0 wbs_dat_o[27]
port 399 nsew signal tristate
flabel metal2 s 194152 -960 194376 480 0 FreeSans 896 90 0 0 wbs_dat_o[28]
port 400 nsew signal tristate
flabel metal2 s 199864 -960 200088 480 0 FreeSans 896 90 0 0 wbs_dat_o[29]
port 401 nsew signal tristate
flabel metal2 s 41832 -960 42056 480 0 FreeSans 896 90 0 0 wbs_dat_o[2]
port 402 nsew signal tristate
flabel metal2 s 205576 -960 205800 480 0 FreeSans 896 90 0 0 wbs_dat_o[30]
port 403 nsew signal tristate
flabel metal2 s 211288 -960 211512 480 0 FreeSans 896 90 0 0 wbs_dat_o[31]
port 404 nsew signal tristate
flabel metal2 s 49448 -960 49672 480 0 FreeSans 896 90 0 0 wbs_dat_o[3]
port 405 nsew signal tristate
flabel metal2 s 57064 -960 57288 480 0 FreeSans 896 90 0 0 wbs_dat_o[4]
port 406 nsew signal tristate
flabel metal2 s 62776 -960 63000 480 0 FreeSans 896 90 0 0 wbs_dat_o[5]
port 407 nsew signal tristate
flabel metal2 s 68488 -960 68712 480 0 FreeSans 896 90 0 0 wbs_dat_o[6]
port 408 nsew signal tristate
flabel metal2 s 74200 -960 74424 480 0 FreeSans 896 90 0 0 wbs_dat_o[7]
port 409 nsew signal tristate
flabel metal2 s 79912 -960 80136 480 0 FreeSans 896 90 0 0 wbs_dat_o[8]
port 410 nsew signal tristate
flabel metal2 s 85624 -960 85848 480 0 FreeSans 896 90 0 0 wbs_dat_o[9]
port 411 nsew signal tristate
flabel metal2 s 28504 -960 28728 480 0 FreeSans 896 90 0 0 wbs_sel_i[0]
port 412 nsew signal input
flabel metal2 s 36120 -960 36344 480 0 FreeSans 896 90 0 0 wbs_sel_i[1]
port 413 nsew signal input
flabel metal2 s 43736 -960 43960 480 0 FreeSans 896 90 0 0 wbs_sel_i[2]
port 414 nsew signal input
flabel metal2 s 51352 -960 51576 480 0 FreeSans 896 90 0 0 wbs_sel_i[3]
port 415 nsew signal input
flabel metal2 s 18984 -960 19208 480 0 FreeSans 896 90 0 0 wbs_stb_i
port 416 nsew signal input
flabel metal2 s 20888 -960 21112 480 0 FreeSans 896 90 0 0 wbs_we_i
port 417 nsew signal input
rlabel via4 565630 580322 565630 580322 0 vdd
rlabel via4 550270 568322 550270 568322 0 vss
rlabel metal3 590562 7112 590562 7112 0 io_in[0]
rlabel metal3 583870 382760 583870 382760 0 io_in[10]
rlabel metal3 593082 443240 593082 443240 0 io_in[11]
rlabel metal3 593138 482888 593138 482888 0 io_in[12]
rlabel metal3 592242 522536 592242 522536 0 io_in[13]
rlabel metal3 584206 554792 584206 554792 0 io_in[14]
rlabel metal2 584696 593082 584696 593082 0 io_in[15]
rlabel metal2 518504 593082 518504 593082 0 io_in[16]
rlabel metal2 452312 593082 452312 593082 0 io_in[17]
rlabel metal2 386120 592242 386120 592242 0 io_in[18]
rlabel metal2 319928 592242 319928 592242 0 io_in[19]
rlabel metal3 593082 46984 593082 46984 0 io_in[1]
rlabel metal2 239176 587230 239176 587230 0 io_in[20]
rlabel metal2 175560 587230 175560 587230 0 io_in[21]
rlabel metal2 121352 592242 121352 592242 0 io_in[22]
rlabel metal3 51744 591304 51744 591304 0 io_in[23]
rlabel metal3 6146 565096 6146 565096 0 io_in[24]
rlabel metal3 6146 522984 6146 522984 0 io_in[25]
rlabel metal3 6146 480872 6146 480872 0 io_in[26]
rlabel metal3 7154 438760 7154 438760 0 io_in[27]
rlabel metal3 7154 396648 7154 396648 0 io_in[28]
rlabel metal3 7154 354536 7154 354536 0 io_in[29]
rlabel metal3 593082 86408 593082 86408 0 io_in[2]
rlabel metal3 6146 312424 6146 312424 0 io_in[30]
rlabel metal3 6146 270312 6146 270312 0 io_in[31]
rlabel metal3 7154 228200 7154 228200 0 io_in[32]
rlabel metal3 7154 186088 7154 186088 0 io_in[33]
rlabel metal3 7154 143976 7154 143976 0 io_in[34]
rlabel metal3 6146 101864 6146 101864 0 io_in[35]
rlabel metal3 2310 79128 2310 79128 0 io_in[36]
rlabel metal3 2254 36904 2254 36904 0 io_in[37]
rlabel metal3 593138 126056 593138 126056 0 io_in[3]
rlabel metal3 583758 146216 583758 146216 0 io_in[4]
rlabel metal3 583814 178472 583814 178472 0 io_in[5]
rlabel metal3 593082 245000 593082 245000 0 io_in[6]
rlabel metal3 590618 284648 590618 284648 0 io_in[7]
rlabel metal3 583814 296744 583814 296744 0 io_in[8]
rlabel metal3 593082 363944 593082 363944 0 io_in[9]
rlabel metal3 592242 33768 592242 33768 0 io_oeb[0]
rlabel metal3 583758 404264 583758 404264 0 io_oeb[10]
rlabel metal3 583758 447272 583758 447272 0 io_oeb[11]
rlabel metal3 583758 490280 583758 490280 0 io_oeb[12]
rlabel metal3 593082 548968 593082 548968 0 io_oeb[13]
rlabel metal3 593082 588616 593082 588616 0 io_oeb[14]
rlabel metal2 525448 587230 525448 587230 0 io_oeb[15]
rlabel metal2 474376 593082 474376 593082 0 io_oeb[16]
rlabel metal2 408296 592242 408296 592242 0 io_oeb[17]
rlabel metal2 334600 588070 334600 588070 0 io_oeb[18]
rlabel metal3 273392 591304 273392 591304 0 io_oeb[19]
rlabel metal4 588952 72072 588952 72072 0 io_oeb[1]
rlabel metal3 208488 591304 208488 591304 0 io_oeb[20]
rlabel metal2 143696 588000 143696 588000 0 io_oeb[21]
rlabel metal3 78792 591304 78792 591304 0 io_oeb[22]
rlabel metal2 11256 592242 11256 592242 0 io_oeb[23]
rlabel metal3 7154 544040 7154 544040 0 io_oeb[24]
rlabel metal3 7154 501928 7154 501928 0 io_oeb[25]
rlabel metal3 3430 474264 3430 474264 0 io_oeb[26]
rlabel metal3 3430 431928 3430 431928 0 io_oeb[27]
rlabel metal3 7266 375592 7266 375592 0 io_oeb[28]
rlabel metal3 7154 333480 7154 333480 0 io_oeb[29]
rlabel metal3 593250 112840 593250 112840 0 io_oeb[2]
rlabel metal3 7154 291368 7154 291368 0 io_oeb[30]
rlabel metal3 3318 262584 3318 262584 0 io_oeb[31]
rlabel metal3 3318 220248 3318 220248 0 io_oeb[32]
rlabel metal3 6202 165032 6202 165032 0 io_oeb[33]
rlabel metal3 6202 122920 6202 122920 0 io_oeb[34]
rlabel metal3 6146 80808 6146 80808 0 io_oeb[35]
rlabel metal3 2758 50904 2758 50904 0 io_oeb[36]
rlabel metal3 3318 8792 3318 8792 0 io_oeb[37]
rlabel metal3 590618 152488 590618 152488 0 io_oeb[3]
rlabel metal3 583870 167720 583870 167720 0 io_oeb[4]
rlabel metal3 583870 199976 583870 199976 0 io_oeb[5]
rlabel metal3 583758 232232 583758 232232 0 io_oeb[6]
rlabel metal3 590562 311080 590562 311080 0 io_oeb[7]
rlabel metal3 583758 318248 583758 318248 0 io_oeb[8]
rlabel metal3 583758 361256 583758 361256 0 io_oeb[9]
rlabel metal3 583758 27944 583758 27944 0 io_out[0]
rlabel metal3 583814 393512 583814 393512 0 io_out[10]
rlabel metal3 590618 456456 590618 456456 0 io_out[11]
rlabel metal3 593082 496104 593082 496104 0 io_out[12]
rlabel metal3 592130 535752 592130 535752 0 io_out[13]
rlabel metal4 591304 570472 591304 570472 0 io_out[14]
rlabel metal2 541352 588126 541352 588126 0 io_out[15]
rlabel metal2 496440 592242 496440 592242 0 io_out[16]
rlabel metal2 430248 592242 430248 592242 0 io_out[17]
rlabel metal2 364056 593082 364056 593082 0 io_out[18]
rlabel metal2 286888 587230 286888 587230 0 io_out[19]
rlabel metal3 588840 60200 588840 60200 0 io_out[1]
rlabel metal2 223272 588070 223272 588070 0 io_out[20]
rlabel metal2 165480 593082 165480 593082 0 io_out[21]
rlabel metal3 97664 591304 97664 591304 0 io_out[22]
rlabel metal2 32704 595672 32704 595672 0 io_out[23]
rlabel metal3 2366 573048 2366 573048 0 io_out[24]
rlabel metal3 6202 512456 6202 512456 0 io_out[25]
rlabel metal3 6202 470344 6202 470344 0 io_out[26]
rlabel metal3 6146 428232 6146 428232 0 io_out[27]
rlabel metal3 6146 386120 6146 386120 0 io_out[28]
rlabel metal3 2310 361368 2310 361368 0 io_out[29]
rlabel metal3 591402 99624 591402 99624 0 io_out[2]
rlabel metal3 6202 301896 6202 301896 0 io_out[30]
rlabel metal3 6202 259784 6202 259784 0 io_out[31]
rlabel metal3 6146 217672 6146 217672 0 io_out[32]
rlabel metal3 6146 175560 6146 175560 0 io_out[33]
rlabel metal3 2310 149688 2310 149688 0 io_out[34]
rlabel metal3 7154 91336 7154 91336 0 io_out[35]
rlabel metal3 2758 65016 2758 65016 0 io_out[36]
rlabel metal3 6146 28168 6146 28168 0 io_out[37]
rlabel metal3 593082 139272 593082 139272 0 io_out[3]
rlabel metal3 583926 156968 583926 156968 0 io_out[4]
rlabel metal3 583758 189224 583758 189224 0 io_out[5]
rlabel metal3 584598 221480 584598 221480 0 io_out[6]
rlabel metal3 593082 297864 593082 297864 0 io_out[7]
rlabel metal3 583870 307496 583870 307496 0 io_out[8]
rlabel metal3 590674 377160 590674 377160 0 io_out[9]
rlabel metal2 213304 2814 213304 2814 0 la_data_in[0]
rlabel metal2 270312 462 270312 462 0 la_data_in[10]
rlabel metal2 276024 2758 276024 2758 0 la_data_in[11]
rlabel metal2 281736 2758 281736 2758 0 la_data_in[12]
rlabel metal2 287448 2198 287448 2198 0 la_data_in[13]
rlabel metal2 293160 2254 293160 2254 0 la_data_in[14]
rlabel metal2 298872 2814 298872 2814 0 la_data_in[15]
rlabel metal2 304584 2254 304584 2254 0 la_data_in[16]
rlabel metal2 310296 2254 310296 2254 0 la_data_in[17]
rlabel metal2 316008 2814 316008 2814 0 la_data_in[18]
rlabel metal2 317352 7042 317352 7042 0 la_data_in[19]
rlabel metal2 219128 462 219128 462 0 la_data_in[1]
rlabel metal2 327432 2198 327432 2198 0 la_data_in[20]
rlabel metal2 333144 3262 333144 3262 0 la_data_in[21]
rlabel metal2 338856 2870 338856 2870 0 la_data_in[22]
rlabel metal2 338856 7042 338856 7042 0 la_data_in[23]
rlabel metal2 350280 2814 350280 2814 0 la_data_in[24]
rlabel metal2 355992 3318 355992 3318 0 la_data_in[25]
rlabel metal2 361704 2814 361704 2814 0 la_data_in[26]
rlabel metal2 360360 7042 360360 7042 0 la_data_in[27]
rlabel metal2 373128 2254 373128 2254 0 la_data_in[28]
rlabel metal2 378840 2310 378840 2310 0 la_data_in[29]
rlabel metal2 224840 2758 224840 2758 0 la_data_in[2]
rlabel metal2 384552 2758 384552 2758 0 la_data_in[30]
rlabel metal2 381864 6370 381864 6370 0 la_data_in[31]
rlabel metal2 387240 6202 387240 6202 0 la_data_in[32]
rlabel metal2 401688 3430 401688 3430 0 la_data_in[33]
rlabel metal2 407400 3262 407400 3262 0 la_data_in[34]
rlabel metal2 403368 6146 403368 6146 0 la_data_in[35]
rlabel metal2 408744 7266 408744 7266 0 la_data_in[36]
rlabel metal2 424536 3206 424536 3206 0 la_data_in[37]
rlabel metal2 430360 3542 430360 3542 0 la_data_in[38]
rlabel metal2 424872 7154 424872 7154 0 la_data_in[39]
rlabel metal2 230552 4270 230552 4270 0 la_data_in[3]
rlabel metal2 430248 6986 430248 6986 0 la_data_in[40]
rlabel metal2 447384 3486 447384 3486 0 la_data_in[41]
rlabel metal2 453096 3206 453096 3206 0 la_data_in[42]
rlabel metal2 446376 7266 446376 7266 0 la_data_in[43]
rlabel metal2 451752 7098 451752 7098 0 la_data_in[44]
rlabel metal2 457128 7378 457128 7378 0 la_data_in[45]
rlabel metal2 475944 3374 475944 3374 0 la_data_in[46]
rlabel metal2 481656 3206 481656 3206 0 la_data_in[47]
rlabel metal2 473256 6426 473256 6426 0 la_data_in[48]
rlabel metal2 478632 6146 478632 6146 0 la_data_in[49]
rlabel metal2 236264 4270 236264 4270 0 la_data_in[4]
rlabel metal2 498792 3150 498792 3150 0 la_data_in[50]
rlabel metal2 504504 2534 504504 2534 0 la_data_in[51]
rlabel metal2 494760 6146 494760 6146 0 la_data_in[52]
rlabel metal2 500136 7266 500136 7266 0 la_data_in[53]
rlabel metal2 505512 7042 505512 7042 0 la_data_in[54]
rlabel metal2 527352 2310 527352 2310 0 la_data_in[55]
rlabel metal2 516264 7378 516264 7378 0 la_data_in[56]
rlabel metal2 521640 7154 521640 7154 0 la_data_in[57]
rlabel metal2 527016 7042 527016 7042 0 la_data_in[58]
rlabel metal2 550200 3486 550200 3486 0 la_data_in[59]
rlabel metal2 241864 2758 241864 2758 0 la_data_in[5]
rlabel metal2 537768 6146 537768 6146 0 la_data_in[60]
rlabel metal2 543144 7210 543144 7210 0 la_data_in[61]
rlabel metal2 548520 7042 548520 7042 0 la_data_in[62]
rlabel metal2 573048 2590 573048 2590 0 la_data_in[63]
rlabel metal2 247464 4256 247464 4256 0 la_data_in[6]
rlabel metal2 253176 4270 253176 4270 0 la_data_in[7]
rlabel metal2 258888 3150 258888 3150 0 la_data_in[8]
rlabel metal2 264600 462 264600 462 0 la_data_in[9]
rlabel metal2 215320 2758 215320 2758 0 la_data_out[0]
rlabel metal2 272216 2758 272216 2758 0 la_data_out[10]
rlabel metal2 277928 2814 277928 2814 0 la_data_out[11]
rlabel metal2 283640 3150 283640 3150 0 la_data_out[12]
rlabel metal2 289352 2254 289352 2254 0 la_data_out[13]
rlabel metal2 292264 6146 292264 6146 0 la_data_out[14]
rlabel metal2 300776 2254 300776 2254 0 la_data_out[15]
rlabel metal2 306488 2310 306488 2310 0 la_data_out[16]
rlabel metal2 312200 2534 312200 2534 0 la_data_out[17]
rlabel metal2 313768 6986 313768 6986 0 la_data_out[18]
rlabel metal2 323624 2758 323624 2758 0 la_data_out[19]
rlabel metal2 221032 462 221032 462 0 la_data_out[1]
rlabel metal2 329336 3206 329336 3206 0 la_data_out[20]
rlabel metal2 335048 2758 335048 2758 0 la_data_out[21]
rlabel metal2 340760 2758 340760 2758 0 la_data_out[22]
rlabel metal2 340648 6986 340648 6986 0 la_data_out[23]
rlabel metal2 352184 2870 352184 2870 0 la_data_out[24]
rlabel metal2 357896 3262 357896 3262 0 la_data_out[25]
rlabel metal2 363608 2870 363608 2870 0 la_data_out[26]
rlabel metal2 362152 6986 362152 6986 0 la_data_out[27]
rlabel metal2 375032 2198 375032 2198 0 la_data_out[28]
rlabel metal2 380744 2422 380744 2422 0 la_data_out[29]
rlabel metal2 226744 2758 226744 2758 0 la_data_out[2]
rlabel metal2 386456 2254 386456 2254 0 la_data_out[30]
rlabel metal2 383656 6314 383656 6314 0 la_data_out[31]
rlabel metal2 397880 2254 397880 2254 0 la_data_out[32]
rlabel metal2 403592 3150 403592 3150 0 la_data_out[33]
rlabel metal2 409304 3206 409304 3206 0 la_data_out[34]
rlabel metal2 405160 6986 405160 6986 0 la_data_out[35]
rlabel metal2 410536 7154 410536 7154 0 la_data_out[36]
rlabel metal2 426440 3150 426440 3150 0 la_data_out[37]
rlabel metal2 432152 3430 432152 3430 0 la_data_out[38]
rlabel metal2 426664 7098 426664 7098 0 la_data_out[39]
rlabel metal2 232456 4270 232456 4270 0 la_data_out[3]
rlabel metal2 432040 7210 432040 7210 0 la_data_out[40]
rlabel metal2 449288 3318 449288 3318 0 la_data_out[41]
rlabel metal2 455000 3150 455000 3150 0 la_data_out[42]
rlabel metal2 448168 6930 448168 6930 0 la_data_out[43]
rlabel metal2 453544 7042 453544 7042 0 la_data_out[44]
rlabel metal2 472136 3486 472136 3486 0 la_data_out[45]
rlabel metal2 477848 3318 477848 3318 0 la_data_out[46]
rlabel metal2 469672 6986 469672 6986 0 la_data_out[47]
rlabel metal2 475048 6314 475048 6314 0 la_data_out[48]
rlabel metal2 480424 6258 480424 6258 0 la_data_out[49]
rlabel metal2 238168 4270 238168 4270 0 la_data_out[4]
rlabel metal2 500696 2646 500696 2646 0 la_data_out[50]
rlabel metal2 491176 6314 491176 6314 0 la_data_out[51]
rlabel metal2 496552 6258 496552 6258 0 la_data_out[52]
rlabel metal2 501928 7154 501928 7154 0 la_data_out[53]
rlabel metal2 523544 3150 523544 3150 0 la_data_out[54]
rlabel metal2 512680 6930 512680 6930 0 la_data_out[55]
rlabel metal2 518056 7266 518056 7266 0 la_data_out[56]
rlabel metal2 523432 7098 523432 7098 0 la_data_out[57]
rlabel metal2 528808 6986 528808 6986 0 la_data_out[58]
rlabel metal2 552216 2646 552216 2646 0 la_data_out[59]
rlabel metal2 243880 4256 243880 4256 0 la_data_out[5]
rlabel metal2 539560 7266 539560 7266 0 la_data_out[60]
rlabel metal2 544936 7154 544936 7154 0 la_data_out[61]
rlabel metal2 550312 6986 550312 6986 0 la_data_out[62]
rlabel metal2 574952 2478 574952 2478 0 la_data_out[63]
rlabel metal2 249368 4270 249368 4270 0 la_data_out[6]
rlabel metal2 255080 4270 255080 4270 0 la_data_out[7]
rlabel metal2 260792 462 260792 462 0 la_data_out[8]
rlabel metal2 266504 2758 266504 2758 0 la_data_out[9]
rlabel metal2 217224 2758 217224 2758 0 la_oenb[0]
rlabel metal2 274120 2758 274120 2758 0 la_oenb[10]
rlabel metal2 279832 2926 279832 2926 0 la_oenb[11]
rlabel metal2 285656 2254 285656 2254 0 la_oenb[12]
rlabel metal2 291256 2198 291256 2198 0 la_oenb[13]
rlabel metal2 296968 2758 296968 2758 0 la_oenb[14]
rlabel metal2 302680 2198 302680 2198 0 la_oenb[15]
rlabel metal2 308392 2422 308392 2422 0 la_oenb[16]
rlabel metal2 314216 2758 314216 2758 0 la_oenb[17]
rlabel metal2 315560 7098 315560 7098 0 la_oenb[18]
rlabel metal2 325528 2254 325528 2254 0 la_oenb[19]
rlabel metal2 222936 3150 222936 3150 0 la_oenb[1]
rlabel metal2 331240 3150 331240 3150 0 la_oenb[20]
rlabel metal2 336952 2814 336952 2814 0 la_oenb[21]
rlabel metal2 337064 7098 337064 7098 0 la_oenb[22]
rlabel metal2 348376 2758 348376 2758 0 la_oenb[23]
rlabel metal2 354088 3150 354088 3150 0 la_oenb[24]
rlabel metal2 359800 2758 359800 2758 0 la_oenb[25]
rlabel metal2 358568 7098 358568 7098 0 la_oenb[26]
rlabel metal2 363944 6258 363944 6258 0 la_oenb[27]
rlabel metal2 376936 2366 376936 2366 0 la_oenb[28]
rlabel metal2 382648 3206 382648 3206 0 la_oenb[29]
rlabel metal2 228648 4270 228648 4270 0 la_oenb[2]
rlabel metal2 380072 6146 380072 6146 0 la_oenb[30]
rlabel metal2 385448 6258 385448 6258 0 la_oenb[31]
rlabel metal2 399896 3374 399896 3374 0 la_oenb[32]
rlabel metal2 405496 3318 405496 3318 0 la_oenb[33]
rlabel metal2 411208 2254 411208 2254 0 la_oenb[34]
rlabel metal2 406952 7210 406952 7210 0 la_oenb[35]
rlabel metal2 422632 2758 422632 2758 0 la_oenb[36]
rlabel metal2 428456 3374 428456 3374 0 la_oenb[37]
rlabel metal2 434056 3486 434056 3486 0 la_oenb[38]
rlabel metal2 429128 7056 429128 7056 0 la_oenb[39]
rlabel metal2 234360 4270 234360 4270 0 la_oenb[3]
rlabel metal2 433832 7266 433832 7266 0 la_oenb[40]
rlabel metal2 451192 3262 451192 3262 0 la_oenb[41]
rlabel metal2 457016 3374 457016 3374 0 la_oenb[42]
rlabel metal2 449960 7154 449960 7154 0 la_oenb[43]
rlabel metal2 455336 6986 455336 6986 0 la_oenb[44]
rlabel metal2 474040 3430 474040 3430 0 la_oenb[45]
rlabel metal2 479752 3262 479752 3262 0 la_oenb[46]
rlabel metal2 471464 6370 471464 6370 0 la_oenb[47]
rlabel metal2 476840 6202 476840 6202 0 la_oenb[48]
rlabel metal2 496888 3206 496888 3206 0 la_oenb[49]
rlabel metal2 240072 2758 240072 2758 0 la_oenb[4]
rlabel metal2 502600 2590 502600 2590 0 la_oenb[50]
rlabel metal2 492968 6202 492968 6202 0 la_oenb[51]
rlabel metal2 498344 7210 498344 7210 0 la_oenb[52]
rlabel metal2 503720 7098 503720 7098 0 la_oenb[53]
rlabel metal2 525448 2366 525448 2366 0 la_oenb[54]
rlabel metal2 514472 7322 514472 7322 0 la_oenb[55]
rlabel metal2 519848 7210 519848 7210 0 la_oenb[56]
rlabel metal2 525224 6370 525224 6370 0 la_oenb[57]
rlabel metal2 548296 2478 548296 2478 0 la_oenb[58]
rlabel metal2 535976 6258 535976 6258 0 la_oenb[59]
rlabel metal2 245672 4256 245672 4256 0 la_oenb[5]
rlabel metal2 541352 6202 541352 6202 0 la_oenb[60]
rlabel metal2 546728 7098 546728 7098 0 la_oenb[61]
rlabel metal2 552104 6370 552104 6370 0 la_oenb[62]
rlabel metal4 557480 5751 557480 5751 0 la_oenb[63]
rlabel metal2 251272 4270 251272 4270 0 la_oenb[6]
rlabel metal2 257096 2758 257096 2758 0 la_oenb[7]
rlabel metal2 262696 462 262696 462 0 la_oenb[8]
rlabel metal2 268408 462 268408 462 0 la_oenb[9]
rlabel metal2 559272 6146 559272 6146 0 user_clock2
rlabel metal4 561064 5605 561064 5605 0 user_irq[0]
rlabel metal2 562856 6258 562856 6258 0 user_irq[1]
rlabel metal2 564648 6202 564648 6202 0 user_irq[2]
rlabel metal2 11592 3150 11592 3150 0 wb_clk_i
rlabel metal2 27048 6146 27048 6146 0 wb_rst_i
rlabel metal2 28840 6202 28840 6202 0 wbs_ack_o
rlabel metal2 23016 2590 23016 2590 0 wbs_adr_i[0]
rlabel metal2 96936 6426 96936 6426 0 wbs_adr_i[10]
rlabel metal2 102312 6202 102312 6202 0 wbs_adr_i[11]
rlabel metal2 99064 2478 99064 2478 0 wbs_adr_i[12]
rlabel metal2 104888 2534 104888 2534 0 wbs_adr_i[13]
rlabel metal2 118440 6146 118440 6146 0 wbs_adr_i[14]
rlabel metal2 123816 6258 123816 6258 0 wbs_adr_i[15]
rlabel metal2 122024 2254 122024 2254 0 wbs_adr_i[16]
rlabel metal2 127624 2422 127624 2422 0 wbs_adr_i[17]
rlabel metal2 133448 2254 133448 2254 0 wbs_adr_i[18]
rlabel metal2 145320 6202 145320 6202 0 wbs_adr_i[19]
rlabel metal2 30632 2310 30632 2310 0 wbs_adr_i[1]
rlabel metal2 144872 2254 144872 2254 0 wbs_adr_i[20]
rlabel metal2 150584 2422 150584 2422 0 wbs_adr_i[21]
rlabel metal2 156184 2198 156184 2198 0 wbs_adr_i[22]
rlabel metal2 166824 6202 166824 6202 0 wbs_adr_i[23]
rlabel metal2 167720 2198 167720 2198 0 wbs_adr_i[24]
rlabel metal2 173432 3206 173432 3206 0 wbs_adr_i[25]
rlabel metal2 179144 2814 179144 2814 0 wbs_adr_i[26]
rlabel metal2 188328 6202 188328 6202 0 wbs_adr_i[27]
rlabel metal2 190568 2814 190568 2814 0 wbs_adr_i[28]
rlabel metal2 196280 2758 196280 2758 0 wbs_adr_i[29]
rlabel metal2 50344 6370 50344 6370 0 wbs_adr_i[2]
rlabel metal2 201992 2758 201992 2758 0 wbs_adr_i[30]
rlabel metal2 207704 2814 207704 2814 0 wbs_adr_i[31]
rlabel metal2 57512 6202 57512 6202 0 wbs_adr_i[3]
rlabel metal2 53480 2590 53480 2590 0 wbs_adr_i[4]
rlabel metal2 59192 2254 59192 2254 0 wbs_adr_i[5]
rlabel metal2 75432 6538 75432 6538 0 wbs_adr_i[6]
rlabel metal2 80808 6202 80808 6202 0 wbs_adr_i[7]
rlabel metal2 76328 2590 76328 2590 0 wbs_adr_i[8]
rlabel metal2 82040 2366 82040 2366 0 wbs_adr_i[9]
rlabel metal2 30632 6258 30632 6258 0 wbs_cyc_i
rlabel metal2 24920 2646 24920 2646 0 wbs_dat_i[0]
rlabel metal2 98728 6370 98728 6370 0 wbs_dat_i[10]
rlabel metal2 95368 2254 95368 2254 0 wbs_dat_i[11]
rlabel metal2 101080 2310 101080 2310 0 wbs_dat_i[12]
rlabel metal2 106792 2198 106792 2198 0 wbs_dat_i[13]
rlabel metal2 120232 6202 120232 6202 0 wbs_dat_i[14]
rlabel metal2 118216 2142 118216 2142 0 wbs_dat_i[15]
rlabel metal2 123928 2534 123928 2534 0 wbs_dat_i[16]
rlabel metal2 129640 2310 129640 2310 0 wbs_dat_i[17]
rlabel metal2 141736 6258 141736 6258 0 wbs_dat_i[18]
rlabel metal2 147112 6314 147112 6314 0 wbs_dat_i[19]
rlabel metal2 32536 2366 32536 2366 0 wbs_dat_i[1]
rlabel metal2 146776 2534 146776 2534 0 wbs_dat_i[20]
rlabel metal2 152488 2310 152488 2310 0 wbs_dat_i[21]
rlabel metal2 158200 2254 158200 2254 0 wbs_dat_i[22]
rlabel metal2 168616 6258 168616 6258 0 wbs_dat_i[23]
rlabel metal2 169624 2254 169624 2254 0 wbs_dat_i[24]
rlabel metal2 175336 3262 175336 3262 0 wbs_dat_i[25]
rlabel metal2 181048 2758 181048 2758 0 wbs_dat_i[26]
rlabel metal2 190120 6986 190120 6986 0 wbs_dat_i[27]
rlabel metal2 192472 2758 192472 2758 0 wbs_dat_i[28]
rlabel metal2 198184 3150 198184 3150 0 wbs_dat_i[29]
rlabel metal2 52136 6426 52136 6426 0 wbs_dat_i[2]
rlabel metal2 203896 2814 203896 2814 0 wbs_dat_i[30]
rlabel metal2 209608 2758 209608 2758 0 wbs_dat_i[31]
rlabel metal2 47768 2422 47768 2422 0 wbs_dat_i[3]
rlabel metal2 55384 2646 55384 2646 0 wbs_dat_i[4]
rlabel metal2 71848 6258 71848 6258 0 wbs_dat_i[5]
rlabel metal2 77224 6370 77224 6370 0 wbs_dat_i[6]
rlabel metal2 72520 2422 72520 2422 0 wbs_dat_i[7]
rlabel metal2 78232 2534 78232 2534 0 wbs_dat_i[8]
rlabel metal2 83944 2254 83944 2254 0 wbs_dat_i[9]
rlabel metal2 26824 2702 26824 2702 0 wbs_dat_o[0]
rlabel metal2 100520 6146 100520 6146 0 wbs_dat_o[10]
rlabel metal2 97272 2422 97272 2422 0 wbs_dat_o[11]
rlabel metal2 102984 2366 102984 2366 0 wbs_dat_o[12]
rlabel metal2 108696 2254 108696 2254 0 wbs_dat_o[13]
rlabel metal2 122024 6370 122024 6370 0 wbs_dat_o[14]
rlabel metal2 120120 2198 120120 2198 0 wbs_dat_o[15]
rlabel metal2 125832 2590 125832 2590 0 wbs_dat_o[16]
rlabel metal2 131544 2198 131544 2198 0 wbs_dat_o[17]
rlabel metal2 143528 6146 143528 6146 0 wbs_dat_o[18]
rlabel metal2 142968 2198 142968 2198 0 wbs_dat_o[19]
rlabel metal2 34440 2422 34440 2422 0 wbs_dat_o[1]
rlabel metal2 148680 2478 148680 2478 0 wbs_dat_o[20]
rlabel metal2 154392 2142 154392 2142 0 wbs_dat_o[21]
rlabel metal2 165032 6146 165032 6146 0 wbs_dat_o[22]
rlabel metal2 165816 2310 165816 2310 0 wbs_dat_o[23]
rlabel metal2 171528 2758 171528 2758 0 wbs_dat_o[24]
rlabel metal2 177240 2870 177240 2870 0 wbs_dat_o[25]
rlabel metal2 182952 2254 182952 2254 0 wbs_dat_o[26]
rlabel metal2 188664 2758 188664 2758 0 wbs_dat_o[27]
rlabel metal2 194376 2814 194376 2814 0 wbs_dat_o[28]
rlabel metal2 200088 2814 200088 2814 0 wbs_dat_o[29]
rlabel metal2 53928 6482 53928 6482 0 wbs_dat_o[2]
rlabel metal2 205800 2758 205800 2758 0 wbs_dat_o[30]
rlabel metal2 213416 7042 213416 7042 0 wbs_dat_o[31]
rlabel metal2 49672 2478 49672 2478 0 wbs_dat_o[3]
rlabel metal2 57288 2310 57288 2310 0 wbs_dat_o[4]
rlabel metal2 73640 6314 73640 6314 0 wbs_dat_o[5]
rlabel metal2 79016 6146 79016 6146 0 wbs_dat_o[6]
rlabel metal2 74424 2478 74424 2478 0 wbs_dat_o[7]
rlabel metal2 80136 2310 80136 2310 0 wbs_dat_o[8]
rlabel metal2 95144 6314 95144 6314 0 wbs_dat_o[9]
rlabel metal2 28728 2254 28728 2254 0 wbs_sel_i[0]
rlabel metal2 48552 6314 48552 6314 0 wbs_sel_i[1]
rlabel metal2 55720 6146 55720 6146 0 wbs_sel_i[2]
rlabel metal2 51576 2534 51576 2534 0 wbs_sel_i[3]
rlabel metal2 32424 6314 32424 6314 0 wbs_stb_i
rlabel metal2 34216 6370 34216 6370 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 596040 596040
<< end >>
